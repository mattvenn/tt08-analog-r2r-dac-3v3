magic
tech sky130A
magscale 1 2
timestamp 1720342921
<< viali >>
rect 4445 18921 4479 18955
rect 6101 18921 6135 18955
rect 949 18785 983 18819
rect 2605 18785 2639 18819
rect 4261 18785 4295 18819
rect 5917 18785 5951 18819
rect 6377 18785 6411 18819
rect 7573 18785 7607 18819
rect 9229 18785 9263 18819
rect 11161 18785 11195 18819
rect 12173 18785 12207 18819
rect 12357 18785 12391 18819
rect 12541 18785 12575 18819
rect 14381 18785 14415 18819
rect 16313 18785 16347 18819
rect 17693 18785 17727 18819
rect 2789 18649 2823 18683
rect 1133 18581 1167 18615
rect 6193 18581 6227 18615
rect 7757 18581 7791 18615
rect 9413 18581 9447 18615
rect 10977 18581 11011 18615
rect 12265 18581 12299 18615
rect 12725 18581 12759 18615
rect 14197 18581 14231 18615
rect 16129 18581 16163 18615
rect 17509 18581 17543 18615
rect 11897 18377 11931 18411
rect 7205 18309 7239 18343
rect 10425 18309 10459 18343
rect 7757 18241 7791 18275
rect 3709 18173 3743 18207
rect 5825 18173 5859 18207
rect 7849 18173 7883 18207
rect 8401 18173 8435 18207
rect 10149 18173 10183 18207
rect 10333 18173 10367 18207
rect 11805 18173 11839 18207
rect 13277 18173 13311 18207
rect 16681 18173 16715 18207
rect 3976 18105 4010 18139
rect 5181 18105 5215 18139
rect 5365 18105 5399 18139
rect 5549 18105 5583 18139
rect 6092 18105 6126 18139
rect 8646 18105 8680 18139
rect 11538 18105 11572 18139
rect 13010 18105 13044 18139
rect 5089 18037 5123 18071
rect 8217 18037 8251 18071
rect 9781 18037 9815 18071
rect 10241 18037 10275 18071
rect 16589 18037 16623 18071
rect 4261 17833 4295 17867
rect 4537 17833 4571 17867
rect 6469 17833 6503 17867
rect 7373 17833 7407 17867
rect 8309 17833 8343 17867
rect 10793 17833 10827 17867
rect 12633 17833 12667 17867
rect 4721 17765 4755 17799
rect 6285 17765 6319 17799
rect 7573 17765 7607 17799
rect 10425 17765 10459 17799
rect 10977 17765 11011 17799
rect 12541 17765 12575 17799
rect 13001 17765 13035 17799
rect 4445 17697 4479 17731
rect 5365 17697 5399 17731
rect 6837 17697 6871 17731
rect 7021 17697 7055 17731
rect 7113 17697 7147 17731
rect 8125 17697 8159 17731
rect 8861 17697 8895 17731
rect 10241 17697 10275 17731
rect 10517 17697 10551 17731
rect 10609 17697 10643 17731
rect 11897 17697 11931 17731
rect 12817 17697 12851 17731
rect 12909 17697 12943 17731
rect 13185 17697 13219 17731
rect 5549 17629 5583 17663
rect 8769 17629 8803 17663
rect 11529 17629 11563 17663
rect 15209 17629 15243 17663
rect 5089 17561 5123 17595
rect 5917 17561 5951 17595
rect 4721 17493 4755 17527
rect 5181 17493 5215 17527
rect 6285 17493 6319 17527
rect 6653 17493 6687 17527
rect 7205 17493 7239 17527
rect 7389 17493 7423 17527
rect 9229 17493 9263 17527
rect 5181 17289 5215 17323
rect 8125 17289 8159 17323
rect 12265 17289 12299 17323
rect 7757 17153 7791 17187
rect 14841 17153 14875 17187
rect 15117 17153 15151 17187
rect 7941 17085 7975 17119
rect 8401 17085 8435 17119
rect 8677 17085 8711 17119
rect 11161 17085 11195 17119
rect 11713 17085 11747 17119
rect 11989 17085 12023 17119
rect 12081 17085 12115 17119
rect 13001 17085 13035 17119
rect 5365 17017 5399 17051
rect 11897 17017 11931 17051
rect 12357 17017 12391 17051
rect 4997 16949 5031 16983
rect 5165 16949 5199 16983
rect 8493 16949 8527 16983
rect 8769 16949 8803 16983
rect 10609 16949 10643 16983
rect 16589 16949 16623 16983
rect 7665 16745 7699 16779
rect 9873 16745 9907 16779
rect 13829 16745 13863 16779
rect 9597 16677 9631 16711
rect 10149 16677 10183 16711
rect 12090 16677 12124 16711
rect 12694 16677 12728 16711
rect 3709 16609 3743 16643
rect 3976 16609 4010 16643
rect 5365 16609 5399 16643
rect 5549 16609 5583 16643
rect 6285 16609 6319 16643
rect 6552 16609 6586 16643
rect 8309 16609 8343 16643
rect 8677 16609 8711 16643
rect 9229 16609 9263 16643
rect 9322 16609 9356 16643
rect 9505 16609 9539 16643
rect 9735 16609 9769 16643
rect 9965 16609 9999 16643
rect 10241 16609 10275 16643
rect 10333 16609 10367 16643
rect 12449 16609 12483 16643
rect 8861 16541 8895 16575
rect 8953 16541 8987 16575
rect 12357 16541 12391 16575
rect 5089 16473 5123 16507
rect 5181 16405 5215 16439
rect 7757 16405 7791 16439
rect 8493 16405 8527 16439
rect 10517 16405 10551 16439
rect 10977 16405 11011 16439
rect 4353 16201 4387 16235
rect 4905 16201 4939 16235
rect 5549 16201 5583 16235
rect 6745 16201 6779 16235
rect 7849 16201 7883 16235
rect 10057 16201 10091 16235
rect 5273 16133 5307 16167
rect 11897 16133 11931 16167
rect 8677 16065 8711 16099
rect 8953 16065 8987 16099
rect 9505 16065 9539 16099
rect 4537 15997 4571 16031
rect 7389 15997 7423 16031
rect 7481 15997 7515 16031
rect 7665 15997 7699 16031
rect 7941 15997 7975 16031
rect 8585 15997 8619 16031
rect 9137 15997 9171 16031
rect 9320 15997 9354 16031
rect 9413 15997 9447 16031
rect 9689 15997 9723 16031
rect 10149 15997 10183 16031
rect 11161 15997 11195 16031
rect 11345 15997 11379 16031
rect 11621 15997 11655 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 13553 15997 13587 16031
rect 13737 15997 13771 16031
rect 5533 15929 5567 15963
rect 5733 15929 5767 15963
rect 11529 15929 11563 15963
rect 12234 15929 12268 15963
rect 4721 15861 4755 15895
rect 4905 15861 4939 15895
rect 5365 15861 5399 15895
rect 9781 15861 9815 15895
rect 10609 15861 10643 15895
rect 13369 15861 13403 15895
rect 13553 15861 13587 15895
rect 10517 15657 10551 15691
rect 10977 15657 11011 15691
rect 12449 15657 12483 15691
rect 5825 15589 5859 15623
rect 6009 15589 6043 15623
rect 7665 15589 7699 15623
rect 7757 15589 7791 15623
rect 8033 15589 8067 15623
rect 10149 15589 10183 15623
rect 12090 15589 12124 15623
rect 2329 15521 2363 15555
rect 2596 15521 2630 15555
rect 4169 15521 4203 15555
rect 7573 15521 7607 15555
rect 7941 15521 7975 15555
rect 9045 15521 9079 15555
rect 9138 15521 9172 15555
rect 9321 15521 9355 15555
rect 9413 15521 9447 15555
rect 9551 15521 9585 15555
rect 9965 15521 9999 15555
rect 10241 15521 10275 15555
rect 10333 15521 10367 15555
rect 13093 15521 13127 15555
rect 4261 15453 4295 15487
rect 8585 15453 8619 15487
rect 12357 15453 12391 15487
rect 3801 15385 3835 15419
rect 3709 15317 3743 15351
rect 6193 15317 6227 15351
rect 7389 15317 7423 15351
rect 9689 15317 9723 15351
rect 2881 15113 2915 15147
rect 6377 15113 6411 15147
rect 6745 14977 6779 15011
rect 3065 14909 3099 14943
rect 3249 14909 3283 14943
rect 3433 14909 3467 14943
rect 3617 14909 3651 14943
rect 4721 14909 4755 14943
rect 4997 14909 5031 14943
rect 7012 14909 7046 14943
rect 8585 14909 8619 14943
rect 11253 14909 11287 14943
rect 11437 14909 11471 14943
rect 11805 14909 11839 14943
rect 11989 14909 12023 14943
rect 13737 14909 13771 14943
rect 13921 14909 13955 14943
rect 5242 14841 5276 14875
rect 8401 14841 8435 14875
rect 11897 14841 11931 14875
rect 4905 14773 4939 14807
rect 8125 14773 8159 14807
rect 8769 14773 8803 14807
rect 11345 14773 11379 14807
rect 13829 14773 13863 14807
rect 3249 14569 3283 14603
rect 3969 14569 4003 14603
rect 5825 14569 5859 14603
rect 7021 14569 7055 14603
rect 11069 14569 11103 14603
rect 13461 14569 13495 14603
rect 3525 14501 3559 14535
rect 4169 14501 4203 14535
rect 6009 14501 6043 14535
rect 7665 14501 7699 14535
rect 8309 14501 8343 14535
rect 8769 14501 8803 14535
rect 1869 14433 1903 14467
rect 2136 14433 2170 14467
rect 3341 14433 3375 14467
rect 6377 14433 6411 14467
rect 6929 14433 6963 14467
rect 7389 14433 7423 14467
rect 7482 14433 7516 14467
rect 7757 14433 7791 14467
rect 7895 14433 7929 14467
rect 8125 14433 8159 14467
rect 8401 14433 8435 14467
rect 8493 14433 8527 14467
rect 9965 14433 9999 14467
rect 10149 14433 10183 14467
rect 10977 14433 11011 14467
rect 11253 14433 11287 14467
rect 11437 14433 11471 14467
rect 11621 14433 11655 14467
rect 13369 14433 13403 14467
rect 13912 14433 13946 14467
rect 9413 14365 9447 14399
rect 13645 14365 13679 14399
rect 15669 14365 15703 14399
rect 3709 14297 3743 14331
rect 8677 14297 8711 14331
rect 15025 14297 15059 14331
rect 3801 14229 3835 14263
rect 3985 14229 4019 14263
rect 6009 14229 6043 14263
rect 8033 14229 8067 14263
rect 10057 14229 10091 14263
rect 11529 14229 11563 14263
rect 15117 14229 15151 14263
rect 2329 14025 2363 14059
rect 3985 14025 4019 14059
rect 4445 14025 4479 14059
rect 5181 14025 5215 14059
rect 7297 14025 7331 14059
rect 7941 14025 7975 14059
rect 8125 14025 8159 14059
rect 10057 14025 10091 14059
rect 13553 14025 13587 14059
rect 14473 14025 14507 14059
rect 3341 13957 3375 13991
rect 8493 13957 8527 13991
rect 11345 13957 11379 13991
rect 4077 13889 4111 13923
rect 12265 13889 12299 13923
rect 13093 13889 13127 13923
rect 13829 13889 13863 13923
rect 2513 13821 2547 13855
rect 3249 13821 3283 13855
rect 3433 13821 3467 13855
rect 3985 13821 4019 13855
rect 4261 13821 4295 13855
rect 7205 13821 7239 13855
rect 7389 13821 7423 13855
rect 7573 13821 7607 13855
rect 7757 13821 7791 13855
rect 8033 13821 8067 13855
rect 8217 13821 8251 13855
rect 8401 13821 8435 13855
rect 8677 13821 8711 13855
rect 11621 13821 11655 13855
rect 12173 13821 12207 13855
rect 13921 13821 13955 13855
rect 14197 13821 14231 13855
rect 14381 13821 14415 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 15025 13821 15059 13855
rect 5135 13787 5169 13821
rect 5365 13753 5399 13787
rect 5917 13753 5951 13787
rect 6101 13753 6135 13787
rect 8944 13753 8978 13787
rect 11345 13753 11379 13787
rect 11529 13753 11563 13787
rect 12081 13753 12115 13787
rect 4997 13685 5031 13719
rect 6285 13685 6319 13719
rect 11713 13685 11747 13719
rect 12541 13685 12575 13719
rect 12909 13685 12943 13719
rect 13001 13685 13035 13719
rect 3065 13481 3099 13515
rect 4629 13481 4663 13515
rect 4905 13481 4939 13515
rect 12265 13481 12299 13515
rect 2697 13413 2731 13447
rect 6561 13413 6595 13447
rect 7297 13413 7331 13447
rect 9045 13413 9079 13447
rect 10977 13413 11011 13447
rect 2421 13345 2455 13379
rect 2605 13345 2639 13379
rect 2881 13345 2915 13379
rect 2973 13345 3007 13379
rect 3249 13345 3283 13379
rect 4261 13345 4295 13379
rect 5089 13345 5123 13379
rect 5181 13345 5215 13379
rect 5365 13345 5399 13379
rect 6193 13345 6227 13379
rect 6837 13345 6871 13379
rect 7021 13345 7055 13379
rect 7205 13345 7239 13379
rect 9229 13345 9263 13379
rect 9597 13345 9631 13379
rect 10149 13345 10183 13379
rect 13461 13345 13495 13379
rect 13645 13345 13679 13379
rect 13737 13345 13771 13379
rect 13829 13345 13863 13379
rect 2697 13277 2731 13311
rect 3433 13277 3467 13311
rect 3525 13277 3559 13311
rect 4169 13277 4203 13311
rect 5273 13277 5307 13311
rect 9689 13277 9723 13311
rect 9873 13277 9907 13311
rect 6745 13209 6779 13243
rect 2421 13141 2455 13175
rect 4629 13141 4663 13175
rect 4813 13141 4847 13175
rect 6561 13141 6595 13175
rect 10333 13141 10367 13175
rect 14105 13141 14139 13175
rect 5181 12937 5215 12971
rect 8217 12937 8251 12971
rect 9689 12937 9723 12971
rect 12173 12937 12207 12971
rect 10333 12869 10367 12903
rect 10701 12869 10735 12903
rect 11805 12869 11839 12903
rect 13093 12869 13127 12903
rect 3801 12801 3835 12835
rect 6837 12801 6871 12835
rect 9873 12801 9907 12835
rect 5549 12733 5583 12767
rect 6009 12733 6043 12767
rect 6653 12733 6687 12767
rect 9597 12733 9631 12767
rect 10060 12733 10094 12767
rect 10333 12733 10367 12767
rect 10593 12711 10627 12745
rect 10701 12733 10735 12767
rect 10885 12733 10919 12767
rect 12081 12733 12115 12767
rect 12357 12733 12391 12767
rect 12449 12733 12483 12767
rect 13093 12733 13127 12767
rect 13369 12733 13403 12767
rect 4068 12665 4102 12699
rect 5917 12665 5951 12699
rect 7104 12665 7138 12699
rect 11805 12665 11839 12699
rect 12173 12665 12207 12699
rect 13277 12665 13311 12699
rect 5825 12597 5859 12631
rect 6101 12597 6135 12631
rect 10241 12597 10275 12631
rect 10517 12597 10551 12631
rect 11989 12597 12023 12631
rect 3617 12393 3651 12427
rect 4261 12393 4295 12427
rect 7205 12393 7239 12427
rect 7297 12393 7331 12427
rect 11161 12393 11195 12427
rect 11345 12393 11379 12427
rect 12173 12393 12207 12427
rect 13001 12393 13035 12427
rect 13829 12393 13863 12427
rect 14289 12393 14323 12427
rect 10333 12325 10367 12359
rect 10517 12325 10551 12359
rect 10977 12325 11011 12359
rect 11805 12325 11839 12359
rect 12633 12325 12667 12359
rect 13461 12325 13495 12359
rect 2237 12257 2271 12291
rect 2504 12257 2538 12291
rect 4445 12257 4479 12291
rect 6081 12257 6115 12291
rect 7481 12257 7515 12291
rect 10609 12257 10643 12291
rect 11253 12257 11287 12291
rect 11713 12257 11747 12291
rect 12541 12257 12575 12291
rect 13369 12257 13403 12291
rect 14197 12257 14231 12291
rect 5825 12189 5859 12223
rect 11897 12189 11931 12223
rect 12725 12189 12759 12223
rect 13553 12189 13587 12223
rect 14381 12189 14415 12223
rect 10333 12053 10367 12087
rect 10977 12053 11011 12087
rect 5733 11849 5767 11883
rect 6101 11849 6135 11883
rect 11621 11849 11655 11883
rect 13185 11849 13219 11883
rect 13553 11849 13587 11883
rect 6837 11713 6871 11747
rect 12265 11713 12299 11747
rect 14381 11713 14415 11747
rect 5917 11645 5951 11679
rect 6193 11645 6227 11679
rect 9321 11645 9355 11679
rect 9505 11645 9539 11679
rect 9689 11645 9723 11679
rect 12081 11645 12115 11679
rect 13921 11645 13955 11679
rect 14013 11645 14047 11679
rect 14197 11645 14231 11679
rect 7082 11577 7116 11611
rect 11989 11577 12023 11611
rect 13001 11577 13035 11611
rect 13737 11577 13771 11611
rect 14105 11577 14139 11611
rect 14626 11577 14660 11611
rect 8217 11509 8251 11543
rect 13206 11509 13240 11543
rect 13369 11509 13403 11543
rect 15761 11509 15795 11543
rect 5273 11305 5307 11339
rect 10057 11305 10091 11339
rect 10701 11305 10735 11339
rect 11897 11305 11931 11339
rect 12265 11305 12299 11339
rect 14013 11305 14047 11339
rect 14565 11305 14599 11339
rect 10425 11237 10459 11271
rect 10517 11237 10551 11271
rect 13645 11237 13679 11271
rect 10195 11203 10229 11237
rect 3893 11169 3927 11203
rect 4149 11169 4183 11203
rect 8493 11169 8527 11203
rect 8760 11169 8794 11203
rect 10793 11169 10827 11203
rect 12081 11169 12115 11203
rect 12357 11169 12391 11203
rect 13461 11169 13495 11203
rect 13737 11169 13771 11203
rect 13829 11169 13863 11203
rect 14381 11169 14415 11203
rect 10517 11033 10551 11067
rect 9873 10965 9907 10999
rect 10241 10965 10275 10999
rect 4077 10761 4111 10795
rect 6929 10761 6963 10795
rect 8861 10761 8895 10795
rect 9505 10761 9539 10795
rect 5549 10693 5583 10727
rect 10149 10693 10183 10727
rect 11069 10693 11103 10727
rect 4537 10625 4571 10659
rect 4997 10625 5031 10659
rect 6377 10625 6411 10659
rect 9597 10625 9631 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 4261 10557 4295 10591
rect 4353 10557 4387 10591
rect 4629 10557 4663 10591
rect 5089 10557 5123 10591
rect 6285 10557 6319 10591
rect 6748 10557 6782 10591
rect 7021 10557 7055 10591
rect 7205 10557 7239 10591
rect 7481 10557 7515 10591
rect 9321 10557 9355 10591
rect 10333 10557 10367 10591
rect 10425 10557 10459 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 10793 10557 10827 10591
rect 10885 10557 10919 10591
rect 11069 10557 11103 10591
rect 11161 10557 11195 10591
rect 15577 10557 15611 10591
rect 16037 10557 16071 10591
rect 7665 10489 7699 10523
rect 8953 10489 8987 10523
rect 9137 10489 9171 10523
rect 5181 10421 5215 10455
rect 6745 10421 6779 10455
rect 11253 10421 11287 10455
rect 15945 10421 15979 10455
rect 16129 10421 16163 10455
rect 3817 10217 3851 10251
rect 3985 10217 4019 10251
rect 6745 10217 6779 10251
rect 7481 10217 7515 10251
rect 7665 10217 7699 10251
rect 11989 10217 12023 10251
rect 13645 10217 13679 10251
rect 16221 10217 16255 10251
rect 3617 10149 3651 10183
rect 15025 10149 15059 10183
rect 4264 10081 4298 10115
rect 4353 10081 4387 10115
rect 4537 10081 4571 10115
rect 4629 10081 4663 10115
rect 5273 10081 5307 10115
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 6285 10081 6319 10115
rect 6561 10081 6595 10115
rect 7113 10081 7147 10115
rect 7849 10081 7883 10115
rect 7941 10081 7975 10115
rect 8125 10081 8159 10115
rect 8217 10081 8251 10115
rect 9137 10081 9171 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 11437 10081 11471 10115
rect 12265 10081 12299 10115
rect 12357 10081 12391 10115
rect 12449 10081 12483 10115
rect 12633 10081 12667 10115
rect 12909 10081 12943 10115
rect 13093 10081 13127 10115
rect 13185 10081 13219 10115
rect 13461 10081 13495 10115
rect 13737 10081 13771 10115
rect 14836 10081 14870 10115
rect 14933 10081 14967 10115
rect 15208 10081 15242 10115
rect 15301 10081 15335 10115
rect 15393 10081 15427 10115
rect 15577 10081 15611 10115
rect 16129 10081 16163 10115
rect 16313 10081 16347 10115
rect 4997 10013 5031 10047
rect 6469 10013 6503 10047
rect 7021 10013 7055 10047
rect 7205 10013 7239 10047
rect 7297 10013 7331 10047
rect 11069 10013 11103 10047
rect 13277 10013 13311 10047
rect 14013 10013 14047 10047
rect 5457 9945 5491 9979
rect 9045 9945 9079 9979
rect 14657 9945 14691 9979
rect 15393 9945 15427 9979
rect 3801 9877 3835 9911
rect 4077 9877 4111 9911
rect 4721 9877 4755 9911
rect 5181 9877 5215 9911
rect 6285 9877 6319 9911
rect 13829 9877 13863 9911
rect 13921 9877 13955 9911
rect 4629 9673 4663 9707
rect 6377 9673 6411 9707
rect 6745 9673 6779 9707
rect 7205 9673 7239 9707
rect 11161 9673 11195 9707
rect 12173 9673 12207 9707
rect 13093 9673 13127 9707
rect 13553 9673 13587 9707
rect 15117 9673 15151 9707
rect 6285 9605 6319 9639
rect 6653 9605 6687 9639
rect 7297 9605 7331 9639
rect 9781 9605 9815 9639
rect 15853 9605 15887 9639
rect 16589 9605 16623 9639
rect 4905 9537 4939 9571
rect 5089 9537 5123 9571
rect 6469 9537 6503 9571
rect 6561 9537 6595 9571
rect 7113 9537 7147 9571
rect 11529 9537 11563 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 4813 9469 4847 9503
rect 4997 9469 5031 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 7389 9469 7423 9503
rect 7481 9469 7515 9503
rect 7665 9469 7699 9503
rect 8953 9469 8987 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 11069 9469 11103 9503
rect 11345 9469 11379 9503
rect 11437 9469 11471 9503
rect 11621 9469 11655 9503
rect 12353 9469 12387 9503
rect 12449 9469 12483 9503
rect 12817 9469 12851 9503
rect 12909 9469 12943 9503
rect 13093 9469 13127 9503
rect 13737 9469 13771 9503
rect 13829 9469 13863 9503
rect 14039 9469 14073 9503
rect 14197 9469 14231 9503
rect 14657 9469 14691 9503
rect 14933 9469 14967 9503
rect 15209 9469 15243 9503
rect 15302 9469 15336 9503
rect 15485 9469 15519 9503
rect 15715 9469 15749 9503
rect 15945 9469 15979 9503
rect 16129 9469 16163 9503
rect 16221 9469 16255 9503
rect 16405 9469 16439 9503
rect 16497 9469 16531 9503
rect 16865 9469 16899 9503
rect 7573 9401 7607 9435
rect 13921 9401 13955 9435
rect 15577 9401 15611 9435
rect 16589 9401 16623 9435
rect 8769 9333 8803 9367
rect 13277 9333 13311 9367
rect 14749 9333 14783 9367
rect 16773 9333 16807 9367
rect 7113 9129 7147 9163
rect 8861 9129 8895 9163
rect 11345 9129 11379 9163
rect 13093 9129 13127 9163
rect 13737 9129 13771 9163
rect 6745 9061 6779 9095
rect 6945 9061 6979 9095
rect 8033 9061 8067 9095
rect 8493 9061 8527 9095
rect 8585 9061 8619 9095
rect 9029 9061 9063 9095
rect 9229 9061 9263 9095
rect 9873 9061 9907 9095
rect 7389 8993 7423 9027
rect 7573 8993 7607 9027
rect 7849 8993 7883 9027
rect 8109 8983 8143 9017
rect 8355 8993 8389 9027
rect 8769 8993 8803 9027
rect 9505 8993 9539 9027
rect 9597 8993 9631 9027
rect 9689 8993 9723 9027
rect 9781 8993 9815 9027
rect 9965 8993 9999 9027
rect 11161 8993 11195 9027
rect 11529 8993 11563 9027
rect 11805 8993 11839 9027
rect 12541 8993 12575 9027
rect 12633 8993 12667 9027
rect 12725 8993 12759 9027
rect 12909 8993 12943 9027
rect 13093 8993 13127 9027
rect 13185 8993 13219 9027
rect 13277 8993 13311 9027
rect 13461 8993 13495 9027
rect 13553 8993 13587 9027
rect 13829 8993 13863 9027
rect 14105 8993 14139 9027
rect 15393 8993 15427 9027
rect 15577 8993 15611 9027
rect 16497 8993 16531 9027
rect 16957 8993 16991 9027
rect 17141 8993 17175 9027
rect 13921 8925 13955 8959
rect 16313 8925 16347 8959
rect 7665 8857 7699 8891
rect 6929 8789 6963 8823
rect 7481 8789 7515 8823
rect 8217 8789 8251 8823
rect 9023 8789 9057 8823
rect 11621 8789 11655 8823
rect 14289 8789 14323 8823
rect 15393 8789 15427 8823
rect 16681 8789 16715 8823
rect 16773 8789 16807 8823
rect 4261 8585 4295 8619
rect 5825 8585 5859 8619
rect 9137 8585 9171 8619
rect 9413 8585 9447 8619
rect 13553 8585 13587 8619
rect 14841 8585 14875 8619
rect 3617 8517 3651 8551
rect 9229 8517 9263 8551
rect 10885 8517 10919 8551
rect 10977 8517 11011 8551
rect 14473 8517 14507 8551
rect 15945 8517 15979 8551
rect 4445 8449 4479 8483
rect 4813 8449 4847 8483
rect 5457 8449 5491 8483
rect 9505 8449 9539 8483
rect 9873 8449 9907 8483
rect 10333 8449 10367 8483
rect 11989 8449 12023 8483
rect 16497 8449 16531 8483
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 4261 8381 4295 8415
rect 4629 8381 4663 8415
rect 4721 8381 4755 8415
rect 4905 8381 4939 8415
rect 5181 8381 5215 8415
rect 5273 8381 5307 8415
rect 5549 8381 5583 8415
rect 6009 8381 6043 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 6377 8381 6411 8415
rect 6561 8381 6595 8415
rect 6929 8381 6963 8415
rect 7205 8381 7239 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 10057 8381 10091 8415
rect 10701 8381 10735 8415
rect 11621 8381 11655 8415
rect 11805 8381 11839 8415
rect 13737 8381 13771 8415
rect 13829 8381 13863 8415
rect 14197 8381 14231 8415
rect 14657 8381 14691 8415
rect 14841 8381 14875 8415
rect 15025 8381 15059 8415
rect 15209 8381 15243 8415
rect 16313 8381 16347 8415
rect 3893 8313 3927 8347
rect 4537 8313 4571 8347
rect 4997 8313 5031 8347
rect 6837 8313 6871 8347
rect 8953 8313 8987 8347
rect 9137 8313 9171 8347
rect 11161 8313 11195 8347
rect 11345 8313 11379 8347
rect 11529 8313 11563 8347
rect 13921 8313 13955 8347
rect 14039 8313 14073 8347
rect 16405 8313 16439 8347
rect 4169 8245 4203 8279
rect 7113 8245 7147 8279
rect 8585 8245 8619 8279
rect 9781 8245 9815 8279
rect 9965 8245 9999 8279
rect 10517 8245 10551 8279
rect 10609 8245 10643 8279
rect 11253 8245 11287 8279
rect 15393 8245 15427 8279
rect 3893 8041 3927 8075
rect 6193 8041 6227 8075
rect 6745 8041 6779 8075
rect 9965 8041 9999 8075
rect 10133 8041 10167 8075
rect 12909 8041 12943 8075
rect 13369 8041 13403 8075
rect 15025 8041 15059 8075
rect 4629 7973 4663 8007
rect 5089 7973 5123 8007
rect 5457 7973 5491 8007
rect 10333 7973 10367 8007
rect 12541 7973 12575 8007
rect 17049 7973 17083 8007
rect 17233 7973 17267 8007
rect 3442 7905 3476 7939
rect 3709 7905 3743 7939
rect 4169 7905 4203 7939
rect 4537 7905 4571 7939
rect 4721 7905 4755 7939
rect 4905 7905 4939 7939
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 6101 7905 6135 7939
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 6561 7905 6595 7939
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 9781 7905 9815 7939
rect 9873 7905 9907 7939
rect 13185 7905 13219 7939
rect 13277 7905 13311 7939
rect 13461 7905 13495 7939
rect 15209 7905 15243 7939
rect 15393 7905 15427 7939
rect 15485 7905 15519 7939
rect 15669 7905 15703 7939
rect 15761 7905 15795 7939
rect 15945 7905 15979 7939
rect 16308 7905 16342 7939
rect 16405 7905 16439 7939
rect 16497 7905 16531 7939
rect 16680 7905 16714 7939
rect 16773 7905 16807 7939
rect 3893 7837 3927 7871
rect 5825 7837 5859 7871
rect 12725 7837 12759 7871
rect 12817 7837 12851 7871
rect 13093 7837 13127 7871
rect 16865 7837 16899 7871
rect 16129 7769 16163 7803
rect 2329 7701 2363 7735
rect 4077 7701 4111 7735
rect 4353 7701 4387 7735
rect 6929 7701 6963 7735
rect 9505 7701 9539 7735
rect 9873 7701 9907 7735
rect 10149 7701 10183 7735
rect 15945 7701 15979 7735
rect 3433 7497 3467 7531
rect 3893 7497 3927 7531
rect 5089 7497 5123 7531
rect 5733 7497 5767 7531
rect 6377 7497 6411 7531
rect 8401 7497 8435 7531
rect 11345 7497 11379 7531
rect 12633 7497 12667 7531
rect 15301 7497 15335 7531
rect 16313 7497 16347 7531
rect 6745 7429 6779 7463
rect 7849 7429 7883 7463
rect 13553 7429 13587 7463
rect 12357 7361 12391 7395
rect 14841 7361 14875 7395
rect 3617 7293 3651 7327
rect 3709 7293 3743 7327
rect 3985 7293 4019 7327
rect 4813 7293 4847 7327
rect 4905 7293 4939 7327
rect 5641 7293 5675 7327
rect 5825 7293 5859 7327
rect 6377 7293 6411 7327
rect 6561 7293 6595 7327
rect 6929 7293 6963 7327
rect 7481 7293 7515 7327
rect 7665 7293 7699 7327
rect 7849 7293 7883 7327
rect 8401 7293 8435 7327
rect 8585 7293 8619 7327
rect 11253 7293 11287 7327
rect 12173 7293 12207 7327
rect 12265 7293 12299 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 12909 7293 12943 7327
rect 13185 7293 13219 7327
rect 13829 7293 13863 7327
rect 14473 7293 14507 7327
rect 16313 7293 16347 7327
rect 16497 7293 16531 7327
rect 16589 7293 16623 7327
rect 16773 7293 16807 7327
rect 13093 7225 13127 7259
rect 13553 7225 13587 7259
rect 14657 7225 14691 7259
rect 15209 7225 15243 7259
rect 16681 7225 16715 7259
rect 13737 7157 13771 7191
rect 5549 6953 5583 6987
rect 11069 6953 11103 6987
rect 12081 6953 12115 6987
rect 12725 6953 12759 6987
rect 4997 6817 5031 6851
rect 5365 6817 5399 6851
rect 5457 6817 5491 6851
rect 7021 6817 7055 6851
rect 7205 6817 7239 6851
rect 7481 6817 7515 6851
rect 7665 6817 7699 6851
rect 8033 6817 8067 6851
rect 8125 6817 8159 6851
rect 8309 6817 8343 6851
rect 8841 6817 8875 6851
rect 10517 6817 10551 6851
rect 11161 6817 11195 6851
rect 11437 6817 11471 6851
rect 11989 6817 12023 6851
rect 12173 6817 12207 6851
rect 12633 6817 12667 6851
rect 12817 6817 12851 6851
rect 13277 6817 13311 6851
rect 13461 6817 13495 6851
rect 15209 6817 15243 6851
rect 16313 6817 16347 6851
rect 16497 6817 16531 6851
rect 5089 6749 5123 6783
rect 7573 6749 7607 6783
rect 8585 6749 8619 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 16129 6749 16163 6783
rect 9965 6681 9999 6715
rect 11621 6681 11655 6715
rect 4813 6613 4847 6647
rect 5181 6613 5215 6647
rect 5273 6613 5307 6647
rect 7389 6613 7423 6647
rect 8493 6613 8527 6647
rect 10701 6613 10735 6647
rect 13461 6613 13495 6647
rect 15025 6613 15059 6647
rect 3985 6409 4019 6443
rect 6009 6409 6043 6443
rect 11621 6409 11655 6443
rect 11805 6409 11839 6443
rect 15669 6409 15703 6443
rect 16313 6409 16347 6443
rect 14657 6341 14691 6375
rect 4537 6273 4571 6307
rect 5917 6273 5951 6307
rect 15577 6273 15611 6307
rect 15945 6273 15979 6307
rect 16589 6273 16623 6307
rect 4905 6205 4939 6239
rect 5089 6205 5123 6239
rect 5181 6205 5215 6239
rect 5273 6205 5307 6239
rect 6009 6205 6043 6239
rect 7481 6205 7515 6239
rect 7757 6205 7791 6239
rect 7941 6205 7975 6239
rect 8033 6205 8067 6239
rect 8401 6205 8435 6239
rect 10241 6205 10275 6239
rect 10497 6205 10531 6239
rect 11713 6205 11747 6239
rect 11897 6205 11931 6239
rect 13553 6205 13587 6239
rect 13737 6205 13771 6239
rect 13829 6205 13863 6239
rect 13921 6205 13955 6239
rect 14565 6205 14599 6239
rect 14749 6205 14783 6239
rect 14841 6205 14875 6239
rect 15209 6205 15243 6239
rect 15853 6205 15887 6239
rect 16037 6205 16071 6239
rect 16129 6205 16163 6239
rect 16497 6205 16531 6239
rect 17049 6205 17083 6239
rect 4353 6137 4387 6171
rect 15393 6137 15427 6171
rect 17233 6137 17267 6171
rect 4445 6069 4479 6103
rect 5549 6069 5583 6103
rect 5641 6069 5675 6103
rect 7297 6069 7331 6103
rect 8125 6069 8159 6103
rect 9689 6069 9723 6103
rect 14197 6069 14231 6103
rect 14381 6069 14415 6103
rect 16957 6069 16991 6103
rect 17417 6069 17451 6103
rect 4261 5865 4295 5899
rect 6929 5865 6963 5899
rect 7021 5865 7055 5899
rect 12817 5865 12851 5899
rect 15025 5865 15059 5899
rect 4813 5797 4847 5831
rect 6101 5797 6135 5831
rect 6193 5797 6227 5831
rect 7481 5797 7515 5831
rect 10977 5797 11011 5831
rect 16865 5797 16899 5831
rect 3148 5729 3182 5763
rect 4537 5729 4571 5763
rect 4629 5729 4663 5763
rect 4905 5729 4939 5763
rect 5089 5729 5123 5763
rect 5181 5729 5215 5763
rect 5457 5729 5491 5763
rect 5825 5729 5859 5763
rect 5973 5729 6007 5763
rect 6331 5729 6365 5763
rect 6837 5729 6871 5763
rect 7297 5729 7331 5763
rect 7389 5729 7423 5763
rect 7573 5729 7607 5763
rect 9321 5729 9355 5763
rect 9669 5729 9703 5763
rect 13001 5729 13035 5763
rect 13093 5729 13127 5763
rect 13185 5729 13219 5763
rect 13369 5729 13403 5763
rect 13829 5729 13863 5763
rect 14013 5729 14047 5763
rect 14197 5729 14231 5763
rect 14381 5729 14415 5763
rect 14933 5729 14967 5763
rect 15117 5729 15151 5763
rect 16129 5729 16163 5763
rect 16221 5729 16255 5763
rect 16405 5729 16439 5763
rect 16497 5729 16531 5763
rect 16773 5729 16807 5763
rect 16957 5729 16991 5763
rect 2881 5661 2915 5695
rect 4813 5661 4847 5695
rect 5273 5661 5307 5695
rect 9413 5661 9447 5695
rect 14289 5661 14323 5695
rect 10793 5593 10827 5627
rect 5641 5525 5675 5559
rect 6469 5525 6503 5559
rect 6561 5525 6595 5559
rect 7205 5525 7239 5559
rect 9229 5525 9263 5559
rect 12265 5525 12299 5559
rect 13921 5525 13955 5559
rect 16681 5525 16715 5559
rect 6193 5321 6227 5355
rect 11069 5321 11103 5355
rect 12909 5321 12943 5355
rect 14289 5321 14323 5355
rect 15485 5321 15519 5355
rect 16313 5321 16347 5355
rect 7757 5253 7791 5287
rect 11437 5253 11471 5287
rect 16129 5253 16163 5287
rect 6285 5185 6319 5219
rect 8677 5185 8711 5219
rect 12633 5185 12667 5219
rect 14565 5185 14599 5219
rect 14933 5185 14967 5219
rect 5822 5117 5856 5151
rect 7481 5117 7515 5151
rect 7665 5117 7699 5151
rect 7941 5117 7975 5151
rect 8217 5117 8251 5151
rect 8585 5117 8619 5151
rect 8769 5117 8803 5151
rect 8861 5117 8895 5151
rect 11253 5117 11287 5151
rect 11345 5117 11379 5151
rect 12449 5117 12483 5151
rect 12541 5117 12575 5151
rect 12725 5117 12759 5151
rect 13001 5117 13035 5151
rect 14197 5117 14231 5151
rect 14473 5117 14507 5151
rect 15209 5117 15243 5151
rect 15577 5117 15611 5151
rect 16313 5117 16347 5151
rect 16497 5117 16531 5151
rect 7573 5049 7607 5083
rect 8125 5049 8159 5083
rect 14841 5049 14875 5083
rect 5641 4981 5675 5015
rect 5825 4981 5859 5015
rect 8401 4981 8435 5015
rect 13093 4981 13127 5015
rect 14105 4981 14139 5015
rect 14657 4981 14691 5015
rect 15025 4981 15059 5015
rect 6285 4777 6319 4811
rect 11069 4777 11103 4811
rect 12449 4777 12483 4811
rect 12725 4777 12759 4811
rect 14841 4777 14875 4811
rect 15117 4709 15151 4743
rect 15669 4709 15703 4743
rect 6101 4641 6135 4675
rect 6285 4641 6319 4675
rect 7205 4641 7239 4675
rect 7297 4641 7331 4675
rect 7573 4641 7607 4675
rect 7757 4641 7791 4675
rect 7849 4641 7883 4675
rect 7941 4641 7975 4675
rect 8033 4641 8067 4675
rect 8401 4641 8435 4675
rect 8493 4641 8527 4675
rect 8677 4641 8711 4675
rect 11253 4641 11287 4675
rect 11437 4641 11471 4675
rect 11713 4641 11747 4675
rect 12265 4641 12299 4675
rect 12725 4641 12759 4675
rect 12909 4641 12943 4675
rect 14197 4641 14231 4675
rect 14381 4641 14415 4675
rect 14565 4641 14599 4675
rect 14749 4641 14783 4675
rect 14979 4641 15013 4675
rect 15209 4641 15243 4675
rect 15392 4641 15426 4675
rect 15485 4641 15519 4675
rect 15577 4641 15611 4675
rect 15761 4641 15795 4675
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 12081 4573 12115 4607
rect 12817 4573 12851 4607
rect 13185 4573 13219 4607
rect 14013 4573 14047 4607
rect 14473 4573 14507 4607
rect 7389 4505 7423 4539
rect 11529 4505 11563 4539
rect 13093 4505 13127 4539
rect 8217 4437 8251 4471
rect 8861 4437 8895 4471
rect 11897 4437 11931 4471
rect 8677 4233 8711 4267
rect 12265 4233 12299 4267
rect 14013 4233 14047 4267
rect 14565 4233 14599 4267
rect 13645 4097 13679 4131
rect 5825 4029 5859 4063
rect 8401 4029 8435 4063
rect 9321 4029 9355 4063
rect 10885 4029 10919 4063
rect 12541 4029 12575 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 13737 4029 13771 4063
rect 14473 4029 14507 4063
rect 14657 4029 14691 4063
rect 6070 3961 6104 3995
rect 9566 3961 9600 3995
rect 11152 3961 11186 3995
rect 12357 3961 12391 3995
rect 7205 3893 7239 3927
rect 8861 3893 8895 3927
rect 10701 3893 10735 3927
rect 9873 3689 9907 3723
rect 12357 3689 12391 3723
rect 8493 3553 8527 3587
rect 8760 3553 8794 3587
rect 9965 3553 9999 3587
rect 10977 3553 11011 3587
rect 11233 3553 11267 3587
rect 10149 3417 10183 3451
rect 7757 2601 7791 2635
rect 12817 2601 12851 2635
rect 8892 2533 8926 2567
rect 13952 2533 13986 2567
rect 9137 2397 9171 2431
rect 14197 2397 14231 2431
rect 10057 1853 10091 1887
rect 10324 1785 10358 1819
rect 11437 1717 11471 1751
rect 2605 1513 2639 1547
rect 11805 1513 11839 1547
rect 14657 1513 14691 1547
rect 17877 1513 17911 1547
rect 12918 1445 12952 1479
rect 13522 1445 13556 1479
rect 16764 1445 16798 1479
rect 3729 1377 3763 1411
rect 2237 1309 2271 1343
rect 3985 1309 4019 1343
rect 13185 1309 13219 1343
rect 13277 1309 13311 1343
rect 16497 1309 16531 1343
rect 13645 833 13679 867
rect 13912 765 13946 799
rect 15025 629 15059 663
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18921 4491 18955
rect 4433 18915 4491 18921
rect 6089 18955 6147 18961
rect 6089 18921 6101 18955
rect 6135 18952 6147 18955
rect 10502 18952 10508 18964
rect 6135 18924 10508 18952
rect 6135 18921 6147 18924
rect 6089 18915 6147 18921
rect 4448 18884 4476 18915
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 8386 18884 8392 18896
rect 4448 18856 8392 18884
rect 8386 18844 8392 18856
rect 8444 18844 8450 18896
rect 842 18776 848 18828
rect 900 18816 906 18828
rect 937 18819 995 18825
rect 937 18816 949 18819
rect 900 18788 949 18816
rect 900 18776 906 18788
rect 937 18785 949 18788
rect 983 18785 995 18819
rect 937 18779 995 18785
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 2593 18819 2651 18825
rect 2593 18816 2605 18819
rect 2556 18788 2605 18816
rect 2556 18776 2562 18788
rect 2593 18785 2605 18788
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4212 18788 4261 18816
rect 4212 18776 4218 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5868 18788 5917 18816
rect 5868 18776 5874 18788
rect 5905 18785 5917 18788
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 6362 18776 6368 18828
rect 6420 18776 6426 18828
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7524 18788 7573 18816
rect 7524 18776 7530 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 9180 18788 9229 18816
rect 9180 18776 9186 18788
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 10836 18788 11161 18816
rect 10836 18776 10842 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 12161 18819 12219 18825
rect 12161 18785 12173 18819
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 12176 18748 12204 18779
rect 10152 18720 12204 18748
rect 12360 18748 12388 18779
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12492 18788 12541 18816
rect 12492 18776 12498 18788
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 12529 18779 12587 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14148 18788 14381 18816
rect 14148 18776 14154 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15804 18788 16313 18816
rect 15804 18776 15810 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17460 18788 17693 18816
rect 17460 18776 17466 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 12360 18720 12756 18748
rect 10152 18692 10180 18720
rect 2777 18683 2835 18689
rect 2777 18649 2789 18683
rect 2823 18680 2835 18683
rect 10134 18680 10140 18692
rect 2823 18652 10140 18680
rect 2823 18649 2835 18652
rect 2777 18643 2835 18649
rect 10134 18640 10140 18652
rect 10192 18640 10198 18692
rect 10410 18680 10416 18692
rect 10244 18652 10416 18680
rect 1121 18615 1179 18621
rect 1121 18581 1133 18615
rect 1167 18612 1179 18615
rect 5902 18612 5908 18624
rect 1167 18584 5908 18612
rect 1167 18581 1179 18584
rect 1121 18575 1179 18581
rect 5902 18572 5908 18584
rect 5960 18572 5966 18624
rect 6178 18572 6184 18624
rect 6236 18572 6242 18624
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 8018 18612 8024 18624
rect 7791 18584 8024 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 9401 18615 9459 18621
rect 9401 18581 9413 18615
rect 9447 18612 9459 18615
rect 10244 18612 10272 18652
rect 10410 18640 10416 18652
rect 10468 18640 10474 18692
rect 12176 18680 12204 18720
rect 12526 18680 12532 18692
rect 12176 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 9447 18584 10272 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10376 18584 10977 18612
rect 10376 18572 10382 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 12728 18621 12756 18720
rect 12253 18615 12311 18621
rect 12253 18612 12265 18615
rect 12032 18584 12265 18612
rect 12032 18572 12038 18584
rect 12253 18581 12265 18584
rect 12299 18581 12311 18615
rect 12253 18575 12311 18581
rect 12713 18615 12771 18621
rect 12713 18581 12725 18615
rect 12759 18612 12771 18615
rect 12802 18612 12808 18624
rect 12759 18584 12808 18612
rect 12759 18581 12771 18584
rect 12713 18575 12771 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 13538 18572 13544 18624
rect 13596 18612 13602 18624
rect 14185 18615 14243 18621
rect 14185 18612 14197 18615
rect 13596 18584 14197 18612
rect 13596 18572 13602 18584
rect 14185 18581 14197 18584
rect 14231 18581 14243 18615
rect 14185 18575 14243 18581
rect 16114 18572 16120 18624
rect 16172 18572 16178 18624
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 16724 18584 17509 18612
rect 16724 18572 16730 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 11882 18408 11888 18420
rect 7852 18380 11888 18408
rect 7193 18343 7251 18349
rect 7193 18309 7205 18343
rect 7239 18309 7251 18343
rect 7193 18303 7251 18309
rect 7208 18272 7236 18303
rect 7374 18272 7380 18284
rect 7208 18244 7380 18272
rect 7374 18232 7380 18244
rect 7432 18272 7438 18284
rect 7745 18275 7803 18281
rect 7745 18272 7757 18275
rect 7432 18244 7757 18272
rect 7432 18232 7438 18244
rect 7745 18241 7757 18244
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 7852 18213 7880 18380
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 10413 18343 10471 18349
rect 10413 18340 10425 18343
rect 9732 18312 10425 18340
rect 9732 18300 9738 18312
rect 10413 18309 10425 18312
rect 10459 18340 10471 18343
rect 10778 18340 10784 18352
rect 10459 18312 10784 18340
rect 10459 18309 10471 18312
rect 10413 18303 10471 18309
rect 10778 18300 10784 18312
rect 10836 18300 10842 18352
rect 3697 18207 3755 18213
rect 3697 18173 3709 18207
rect 3743 18204 3755 18207
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 3743 18176 5825 18204
rect 3743 18173 3755 18176
rect 3697 18167 3755 18173
rect 5813 18173 5825 18176
rect 5859 18204 5871 18207
rect 7837 18207 7895 18213
rect 5859 18176 6224 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 3964 18139 4022 18145
rect 3964 18105 3976 18139
rect 4010 18136 4022 18139
rect 4246 18136 4252 18148
rect 4010 18108 4252 18136
rect 4010 18105 4022 18108
rect 3964 18099 4022 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 4706 18096 4712 18148
rect 4764 18136 4770 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 4764 18108 5181 18136
rect 4764 18096 4770 18108
rect 5169 18105 5181 18108
rect 5215 18105 5227 18139
rect 5169 18099 5227 18105
rect 5353 18139 5411 18145
rect 5353 18105 5365 18139
rect 5399 18136 5411 18139
rect 5442 18136 5448 18148
rect 5399 18108 5448 18136
rect 5399 18105 5411 18108
rect 5353 18099 5411 18105
rect 5077 18071 5135 18077
rect 5077 18037 5089 18071
rect 5123 18068 5135 18071
rect 5368 18068 5396 18099
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 5537 18139 5595 18145
rect 5537 18105 5549 18139
rect 5583 18136 5595 18139
rect 5626 18136 5632 18148
rect 5583 18108 5632 18136
rect 5583 18105 5595 18108
rect 5537 18099 5595 18105
rect 5626 18096 5632 18108
rect 5684 18096 5690 18148
rect 6086 18145 6092 18148
rect 6080 18136 6092 18145
rect 6047 18108 6092 18136
rect 6080 18099 6092 18108
rect 6086 18096 6092 18099
rect 6144 18096 6150 18148
rect 6196 18136 6224 18176
rect 7837 18173 7849 18207
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18173 8447 18207
rect 8389 18167 8447 18173
rect 6270 18136 6276 18148
rect 6196 18108 6276 18136
rect 6270 18096 6276 18108
rect 6328 18136 6334 18148
rect 8404 18136 8432 18167
rect 10134 18164 10140 18216
rect 10192 18164 10198 18216
rect 10318 18164 10324 18216
rect 10376 18164 10382 18216
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18204 11851 18207
rect 12066 18204 12072 18216
rect 11839 18176 12072 18204
rect 11839 18173 11851 18176
rect 11793 18167 11851 18173
rect 12066 18164 12072 18176
rect 12124 18204 12130 18216
rect 13265 18207 13323 18213
rect 13265 18204 13277 18207
rect 12124 18176 13277 18204
rect 12124 18164 12130 18176
rect 13265 18173 13277 18176
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 16666 18164 16672 18216
rect 16724 18164 16730 18216
rect 6328 18108 8432 18136
rect 6328 18096 6334 18108
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 8634 18139 8692 18145
rect 8634 18136 8646 18139
rect 8536 18108 8646 18136
rect 8536 18096 8542 18108
rect 8634 18105 8646 18108
rect 8680 18105 8692 18139
rect 8634 18099 8692 18105
rect 11054 18096 11060 18148
rect 11112 18136 11118 18148
rect 11526 18139 11584 18145
rect 11526 18136 11538 18139
rect 11112 18108 11538 18136
rect 11112 18096 11118 18108
rect 11526 18105 11538 18108
rect 11572 18105 11584 18139
rect 11526 18099 11584 18105
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 12998 18139 13056 18145
rect 12998 18136 13010 18139
rect 12676 18108 13010 18136
rect 12676 18096 12682 18108
rect 12998 18105 13010 18108
rect 13044 18105 13056 18139
rect 12998 18099 13056 18105
rect 5123 18040 5396 18068
rect 5123 18037 5135 18040
rect 5077 18031 5135 18037
rect 8202 18028 8208 18080
rect 8260 18028 8266 18080
rect 9582 18028 9588 18080
rect 9640 18068 9646 18080
rect 9769 18071 9827 18077
rect 9769 18068 9781 18071
rect 9640 18040 9781 18068
rect 9640 18028 9646 18040
rect 9769 18037 9781 18040
rect 9815 18037 9827 18071
rect 9769 18031 9827 18037
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 16574 18028 16580 18080
rect 16632 18028 16638 18080
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 4246 17824 4252 17876
rect 4304 17824 4310 17876
rect 4525 17867 4583 17873
rect 4525 17833 4537 17867
rect 4571 17833 4583 17867
rect 4525 17827 4583 17833
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4540 17728 4568 17827
rect 6362 17824 6368 17876
rect 6420 17864 6426 17876
rect 7374 17873 7380 17876
rect 6457 17867 6515 17873
rect 6457 17864 6469 17867
rect 6420 17836 6469 17864
rect 6420 17824 6426 17836
rect 6457 17833 6469 17836
rect 6503 17833 6515 17867
rect 7361 17867 7380 17873
rect 7361 17864 7373 17867
rect 6457 17827 6515 17833
rect 6840 17836 7373 17864
rect 4709 17799 4767 17805
rect 4709 17765 4721 17799
rect 4755 17796 4767 17799
rect 4798 17796 4804 17808
rect 4755 17768 4804 17796
rect 4755 17765 4767 17768
rect 4709 17759 4767 17765
rect 4798 17756 4804 17768
rect 4856 17796 4862 17808
rect 6273 17799 6331 17805
rect 6273 17796 6285 17799
rect 4856 17768 6285 17796
rect 4856 17756 4862 17768
rect 6273 17765 6285 17768
rect 6319 17765 6331 17799
rect 6273 17759 6331 17765
rect 6840 17737 6868 17836
rect 7361 17833 7373 17836
rect 7361 17827 7380 17833
rect 7374 17824 7380 17827
rect 7432 17824 7438 17876
rect 8297 17867 8355 17873
rect 8297 17833 8309 17867
rect 8343 17864 8355 17867
rect 8478 17864 8484 17876
rect 8343 17836 8484 17864
rect 8343 17833 8355 17836
rect 8297 17827 8355 17833
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 10594 17864 10600 17876
rect 10336 17836 10600 17864
rect 7561 17799 7619 17805
rect 6932 17768 7236 17796
rect 4479 17700 4568 17728
rect 5353 17731 5411 17737
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 5353 17697 5365 17731
rect 5399 17697 5411 17731
rect 5353 17691 5411 17697
rect 6825 17731 6883 17737
rect 6825 17697 6837 17731
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17592 5135 17595
rect 5368 17592 5396 17691
rect 5442 17620 5448 17672
rect 5500 17660 5506 17672
rect 5537 17663 5595 17669
rect 5537 17660 5549 17663
rect 5500 17632 5549 17660
rect 5500 17620 5506 17632
rect 5537 17629 5549 17632
rect 5583 17660 5595 17663
rect 6932 17660 6960 17768
rect 7006 17688 7012 17740
rect 7064 17688 7070 17740
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17697 7159 17731
rect 7101 17691 7159 17697
rect 5583 17632 6960 17660
rect 5583 17629 5595 17632
rect 5537 17623 5595 17629
rect 5626 17592 5632 17604
rect 5123 17564 5212 17592
rect 5368 17564 5632 17592
rect 5123 17561 5135 17564
rect 5077 17555 5135 17561
rect 4706 17484 4712 17536
rect 4764 17484 4770 17536
rect 5184 17533 5212 17564
rect 5626 17552 5632 17564
rect 5684 17592 5690 17604
rect 5905 17595 5963 17601
rect 5905 17592 5917 17595
rect 5684 17564 5917 17592
rect 5684 17552 5690 17564
rect 5905 17561 5917 17564
rect 5951 17592 5963 17595
rect 7116 17592 7144 17691
rect 7208 17660 7236 17768
rect 7561 17765 7573 17799
rect 7607 17796 7619 17799
rect 7834 17796 7840 17808
rect 7607 17768 7840 17796
rect 7607 17765 7619 17768
rect 7561 17759 7619 17765
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 8110 17688 8116 17740
rect 8168 17688 8174 17740
rect 8849 17731 8907 17737
rect 8849 17697 8861 17731
rect 8895 17728 8907 17731
rect 9674 17728 9680 17740
rect 8895 17700 9680 17728
rect 8895 17697 8907 17700
rect 8849 17691 8907 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 10229 17731 10287 17737
rect 10229 17697 10241 17731
rect 10275 17697 10287 17731
rect 10336 17728 10364 17836
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 10781 17867 10839 17873
rect 10781 17833 10793 17867
rect 10827 17864 10839 17867
rect 11054 17864 11060 17876
rect 10827 17836 11060 17864
rect 10827 17833 10839 17836
rect 10781 17827 10839 17833
rect 11054 17824 11060 17836
rect 11112 17824 11118 17876
rect 12618 17824 12624 17876
rect 12676 17824 12682 17876
rect 10413 17799 10471 17805
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 10965 17799 11023 17805
rect 10965 17796 10977 17799
rect 10459 17768 10977 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 10965 17765 10977 17768
rect 11011 17765 11023 17799
rect 10965 17759 11023 17765
rect 12529 17799 12587 17805
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12575 17768 13001 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 12989 17765 13001 17768
rect 13035 17765 13047 17799
rect 12989 17759 13047 17765
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 10336 17700 10517 17728
rect 10229 17691 10287 17697
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 10597 17731 10655 17737
rect 10597 17697 10609 17731
rect 10643 17697 10655 17731
rect 10597 17691 10655 17697
rect 8757 17663 8815 17669
rect 8757 17660 8769 17663
rect 7208 17632 8769 17660
rect 8757 17629 8769 17632
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 10244 17592 10272 17691
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10612 17660 10640 17691
rect 11882 17688 11888 17740
rect 11940 17688 11946 17740
rect 12802 17688 12808 17740
rect 12860 17688 12866 17740
rect 12894 17688 12900 17740
rect 12952 17688 12958 17740
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17697 13231 17731
rect 13173 17691 13231 17697
rect 10376 17632 10640 17660
rect 10376 17620 10382 17632
rect 10778 17620 10784 17672
rect 10836 17660 10842 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 10836 17632 11529 17660
rect 10836 17620 10842 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 13188 17660 13216 17691
rect 11517 17623 11575 17629
rect 12406 17632 13216 17660
rect 11054 17592 11060 17604
rect 5951 17564 6776 17592
rect 7116 17564 7420 17592
rect 10244 17564 11060 17592
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 5169 17527 5227 17533
rect 5169 17493 5181 17527
rect 5215 17524 5227 17527
rect 5534 17524 5540 17536
rect 5215 17496 5540 17524
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 6273 17527 6331 17533
rect 6273 17493 6285 17527
rect 6319 17524 6331 17527
rect 6641 17527 6699 17533
rect 6641 17524 6653 17527
rect 6319 17496 6653 17524
rect 6319 17493 6331 17496
rect 6273 17487 6331 17493
rect 6641 17493 6653 17496
rect 6687 17493 6699 17527
rect 6748 17524 6776 17564
rect 7392 17536 7420 17564
rect 11054 17552 11060 17564
rect 11112 17592 11118 17604
rect 12406 17592 12434 17632
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15197 17663 15255 17669
rect 15197 17660 15209 17663
rect 15160 17632 15209 17660
rect 15160 17620 15166 17632
rect 15197 17629 15209 17632
rect 15243 17629 15255 17663
rect 15197 17623 15255 17629
rect 11112 17564 12434 17592
rect 11112 17552 11118 17564
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 6748 17496 7205 17524
rect 6641 17487 6699 17493
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 7374 17484 7380 17536
rect 7432 17484 7438 17536
rect 9214 17484 9220 17536
rect 9272 17484 9278 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5718 17320 5724 17332
rect 5215 17292 5724 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 8110 17280 8116 17332
rect 8168 17280 8174 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12342 17320 12348 17332
rect 12299 17292 12348 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 7006 17212 7012 17264
rect 7064 17252 7070 17264
rect 7834 17252 7840 17264
rect 7064 17224 7840 17252
rect 7064 17212 7070 17224
rect 7834 17212 7840 17224
rect 7892 17252 7898 17264
rect 9674 17252 9680 17264
rect 7892 17224 9680 17252
rect 7892 17212 7898 17224
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 7791 17156 8616 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 4798 17076 4804 17128
rect 4856 17116 4862 17128
rect 7929 17119 7987 17125
rect 7929 17116 7941 17119
rect 4856 17088 7941 17116
rect 4856 17076 4862 17088
rect 7929 17085 7941 17088
rect 7975 17116 7987 17119
rect 8110 17116 8116 17128
rect 7975 17088 8116 17116
rect 7975 17085 7987 17088
rect 7929 17079 7987 17085
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 5353 17051 5411 17057
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 5442 17048 5448 17060
rect 5399 17020 5448 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 8404 17048 8432 17079
rect 7432 17020 8432 17048
rect 8588 17048 8616 17156
rect 8680 17125 8708 17224
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 12894 17252 12900 17264
rect 11992 17224 12900 17252
rect 10226 17144 10232 17196
rect 10284 17184 10290 17196
rect 10594 17184 10600 17196
rect 10284 17156 10600 17184
rect 10284 17144 10290 17156
rect 10594 17144 10600 17156
rect 10652 17184 10658 17196
rect 11606 17184 11612 17196
rect 10652 17156 11612 17184
rect 10652 17144 10658 17156
rect 11606 17144 11612 17156
rect 11664 17184 11670 17196
rect 11992 17184 12020 17224
rect 12894 17212 12900 17224
rect 12952 17212 12958 17264
rect 11664 17156 12020 17184
rect 11664 17144 11670 17156
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17085 8723 17119
rect 8665 17079 8723 17085
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 11992 17125 12020 17156
rect 12250 17144 12256 17196
rect 12308 17184 12314 17196
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 12308 17156 14841 17184
rect 12308 17144 12314 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 11149 17119 11207 17125
rect 11149 17116 11161 17119
rect 11020 17088 11161 17116
rect 11020 17076 11026 17088
rect 11149 17085 11161 17088
rect 11195 17085 11207 17119
rect 11149 17079 11207 17085
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 11977 17119 12035 17125
rect 11977 17085 11989 17119
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12069 17119 12127 17125
rect 12069 17085 12081 17119
rect 12115 17116 12127 17119
rect 12115 17088 12940 17116
rect 12115 17085 12127 17088
rect 12069 17079 12127 17085
rect 8588 17020 8800 17048
rect 7432 17008 7438 17020
rect 4982 16940 4988 16992
rect 5040 16940 5046 16992
rect 5153 16983 5211 16989
rect 5153 16949 5165 16983
rect 5199 16980 5211 16983
rect 5626 16980 5632 16992
rect 5199 16952 5632 16980
rect 5199 16949 5211 16952
rect 5153 16943 5211 16949
rect 5626 16940 5632 16952
rect 5684 16940 5690 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 8772 16989 8800 17020
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 11716 17048 11744 17079
rect 11112 17020 11744 17048
rect 11885 17051 11943 17057
rect 11112 17008 11118 17020
rect 11885 17017 11897 17051
rect 11931 17017 11943 17051
rect 12345 17051 12403 17057
rect 12345 17048 12357 17051
rect 11885 17011 11943 17017
rect 12084 17020 12357 17048
rect 8757 16983 8815 16989
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 9122 16980 9128 16992
rect 8803 16952 9128 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 9122 16940 9128 16952
rect 9180 16940 9186 16992
rect 10410 16940 10416 16992
rect 10468 16980 10474 16992
rect 10597 16983 10655 16989
rect 10597 16980 10609 16983
rect 10468 16952 10609 16980
rect 10468 16940 10474 16952
rect 10597 16949 10609 16952
rect 10643 16949 10655 16983
rect 11900 16980 11928 17011
rect 12084 16980 12112 17020
rect 12345 17017 12357 17020
rect 12391 17017 12403 17051
rect 12912 17048 12940 17088
rect 12986 17076 12992 17128
rect 13044 17076 13050 17128
rect 16574 17116 16580 17128
rect 16238 17088 16580 17116
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 13538 17048 13544 17060
rect 12912 17020 13544 17048
rect 12345 17011 12403 17017
rect 13538 17008 13544 17020
rect 13596 17008 13602 17060
rect 11900 16952 12112 16980
rect 10597 16943 10655 16949
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 16577 16983 16635 16989
rect 16577 16980 16589 16983
rect 12676 16952 16589 16980
rect 12676 16940 12682 16952
rect 16577 16949 16589 16952
rect 16623 16949 16635 16983
rect 16577 16943 16635 16949
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 7653 16779 7711 16785
rect 7653 16776 7665 16779
rect 7432 16748 7665 16776
rect 7432 16736 7438 16748
rect 7653 16745 7665 16748
rect 7699 16745 7711 16779
rect 9674 16776 9680 16788
rect 7653 16739 7711 16745
rect 9600 16748 9680 16776
rect 3712 16680 6316 16708
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 3712 16649 3740 16680
rect 6288 16652 6316 16680
rect 3697 16643 3755 16649
rect 3697 16640 3709 16643
rect 2372 16612 3709 16640
rect 2372 16600 2378 16612
rect 3697 16609 3709 16612
rect 3743 16609 3755 16643
rect 3697 16603 3755 16609
rect 3964 16643 4022 16649
rect 3964 16609 3976 16643
rect 4010 16640 4022 16643
rect 4338 16640 4344 16652
rect 4010 16612 4344 16640
rect 4010 16609 4022 16612
rect 3964 16603 4022 16609
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 5353 16643 5411 16649
rect 5353 16640 5365 16643
rect 5092 16612 5365 16640
rect 5092 16513 5120 16612
rect 5353 16609 5365 16612
rect 5399 16640 5411 16643
rect 5399 16612 5488 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5460 16572 5488 16612
rect 5534 16600 5540 16652
rect 5592 16600 5598 16652
rect 6270 16600 6276 16652
rect 6328 16600 6334 16652
rect 6546 16649 6552 16652
rect 6540 16603 6552 16649
rect 6546 16600 6552 16603
rect 6604 16600 6610 16652
rect 7668 16640 7696 16739
rect 8110 16668 8116 16720
rect 8168 16708 8174 16720
rect 9600 16717 9628 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9861 16779 9919 16785
rect 9861 16745 9873 16779
rect 9907 16776 9919 16779
rect 10594 16776 10600 16788
rect 9907 16748 10600 16776
rect 9907 16745 9919 16748
rect 9861 16739 9919 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 12986 16776 12992 16788
rect 12176 16748 12992 16776
rect 9585 16711 9643 16717
rect 8168 16680 8708 16708
rect 8168 16668 8174 16680
rect 8680 16649 8708 16680
rect 9585 16677 9597 16711
rect 9631 16677 9643 16711
rect 9585 16671 9643 16677
rect 10137 16711 10195 16717
rect 10137 16677 10149 16711
rect 10183 16708 10195 16711
rect 10410 16708 10416 16720
rect 10183 16680 10416 16708
rect 10183 16677 10195 16680
rect 10137 16671 10195 16677
rect 10410 16668 10416 16680
rect 10468 16668 10474 16720
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 12078 16711 12136 16717
rect 12078 16708 12090 16711
rect 10744 16680 12090 16708
rect 10744 16668 10750 16680
rect 12078 16677 12090 16680
rect 12124 16677 12136 16711
rect 12078 16671 12136 16677
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 7668 16612 8309 16640
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 8297 16603 8355 16609
rect 8665 16643 8723 16649
rect 8665 16609 8677 16643
rect 8711 16609 8723 16643
rect 8665 16603 8723 16609
rect 9214 16600 9220 16652
rect 9272 16600 9278 16652
rect 9310 16643 9368 16649
rect 9310 16609 9322 16643
rect 9356 16609 9368 16643
rect 9310 16603 9368 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9723 16643 9781 16649
rect 9539 16612 9628 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 5718 16572 5724 16584
rect 5460 16544 5724 16572
rect 5718 16532 5724 16544
rect 5776 16532 5782 16584
rect 8478 16532 8484 16584
rect 8536 16572 8542 16584
rect 8849 16575 8907 16581
rect 8849 16572 8861 16575
rect 8536 16544 8861 16572
rect 8536 16532 8542 16544
rect 8849 16541 8861 16544
rect 8895 16541 8907 16575
rect 8849 16535 8907 16541
rect 8941 16575 8999 16581
rect 8941 16541 8953 16575
rect 8987 16572 8999 16575
rect 9122 16572 9128 16584
rect 8987 16544 9128 16572
rect 8987 16541 8999 16544
rect 8941 16535 8999 16541
rect 5077 16507 5135 16513
rect 5077 16473 5089 16507
rect 5123 16473 5135 16507
rect 5077 16467 5135 16473
rect 8110 16464 8116 16516
rect 8168 16504 8174 16516
rect 8864 16504 8892 16535
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9324 16504 9352 16603
rect 9600 16572 9628 16612
rect 9723 16609 9735 16643
rect 9769 16640 9781 16643
rect 9858 16640 9864 16652
rect 9769 16612 9864 16640
rect 9769 16609 9781 16612
rect 9723 16603 9781 16609
rect 9858 16600 9864 16612
rect 9916 16600 9922 16652
rect 9950 16600 9956 16652
rect 10008 16600 10014 16652
rect 10226 16600 10232 16652
rect 10284 16600 10290 16652
rect 10318 16600 10324 16652
rect 10376 16600 10382 16652
rect 12176 16640 12204 16748
rect 12986 16736 12992 16748
rect 13044 16776 13050 16788
rect 13817 16779 13875 16785
rect 13817 16776 13829 16779
rect 13044 16748 13829 16776
rect 13044 16736 13050 16748
rect 13817 16745 13829 16748
rect 13863 16745 13875 16779
rect 13817 16739 13875 16745
rect 12342 16668 12348 16720
rect 12400 16708 12406 16720
rect 12682 16711 12740 16717
rect 12682 16708 12694 16711
rect 12400 16680 12694 16708
rect 12400 16668 12406 16680
rect 12682 16677 12694 16680
rect 12728 16677 12740 16711
rect 12682 16671 12740 16677
rect 10428 16612 12204 16640
rect 10428 16572 10456 16612
rect 12250 16600 12256 16652
rect 12308 16640 12314 16652
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 12308 16612 12449 16640
rect 12308 16600 12314 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 9600 16544 10456 16572
rect 12345 16575 12403 16581
rect 9692 16516 9720 16544
rect 12345 16541 12357 16575
rect 12391 16572 12403 16575
rect 12452 16572 12480 16603
rect 12391 16544 12480 16572
rect 12391 16541 12403 16544
rect 12345 16535 12403 16541
rect 9490 16504 9496 16516
rect 8168 16476 8800 16504
rect 8864 16476 9496 16504
rect 8168 16464 8174 16476
rect 5166 16396 5172 16448
rect 5224 16396 5230 16448
rect 7745 16439 7803 16445
rect 7745 16405 7757 16439
rect 7791 16436 7803 16439
rect 7834 16436 7840 16448
rect 7791 16408 7840 16436
rect 7791 16405 7803 16408
rect 7745 16399 7803 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8478 16396 8484 16448
rect 8536 16396 8542 16448
rect 8772 16436 8800 16476
rect 9490 16464 9496 16476
rect 9548 16464 9554 16516
rect 9674 16464 9680 16516
rect 9732 16464 9738 16516
rect 11054 16504 11060 16516
rect 9968 16476 11060 16504
rect 9968 16448 9996 16476
rect 11054 16464 11060 16476
rect 11112 16464 11118 16516
rect 9950 16436 9956 16448
rect 8772 16408 9956 16436
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10505 16439 10563 16445
rect 10505 16405 10517 16439
rect 10551 16436 10563 16439
rect 10686 16436 10692 16448
rect 10551 16408 10692 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 10962 16396 10968 16448
rect 11020 16396 11026 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 12360 16436 12388 16535
rect 12124 16408 12388 16436
rect 12124 16396 12130 16408
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 4338 16192 4344 16244
rect 4396 16192 4402 16244
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5166 16232 5172 16244
rect 4939 16204 5172 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 5537 16235 5595 16241
rect 5537 16201 5549 16235
rect 5583 16232 5595 16235
rect 5994 16232 6000 16244
rect 5583 16204 6000 16232
rect 5583 16201 5595 16204
rect 5537 16195 5595 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 6546 16192 6552 16244
rect 6604 16232 6610 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 6604 16204 6745 16232
rect 6604 16192 6610 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 6733 16195 6791 16201
rect 7834 16192 7840 16244
rect 7892 16192 7898 16244
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 9916 16204 10057 16232
rect 9916 16192 9922 16204
rect 10045 16201 10057 16204
rect 10091 16201 10103 16235
rect 16114 16232 16120 16244
rect 10045 16195 10103 16201
rect 11716 16204 16120 16232
rect 4982 16124 4988 16176
rect 5040 16164 5046 16176
rect 5261 16167 5319 16173
rect 5261 16164 5273 16167
rect 5040 16136 5273 16164
rect 5040 16124 5046 16136
rect 5261 16133 5273 16136
rect 5307 16133 5319 16167
rect 10962 16164 10968 16176
rect 5261 16127 5319 16133
rect 8588 16136 10968 16164
rect 8478 16096 8484 16108
rect 7668 16068 8484 16096
rect 7668 16037 7696 16068
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 7377 16031 7435 16037
rect 4571 16000 4752 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4724 15901 4752 16000
rect 7377 15997 7389 16031
rect 7423 16028 7435 16031
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 7423 16000 7481 16028
rect 7423 15997 7435 16000
rect 7377 15991 7435 15997
rect 7469 15997 7481 16000
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8588 16037 8616 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11112 16136 11376 16164
rect 11112 16124 11118 16136
rect 8662 16056 8668 16108
rect 8720 16056 8726 16108
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9030 16096 9036 16108
rect 8987 16068 9036 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 9640 16068 11284 16096
rect 9640 16056 9646 16068
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 15997 8631 16031
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8573 15991 8631 15997
rect 8680 16000 9137 16028
rect 5534 15969 5540 15972
rect 5521 15963 5540 15969
rect 5521 15929 5533 15963
rect 5521 15923 5540 15929
rect 5534 15920 5540 15923
rect 5592 15920 5598 15972
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 5776 15932 6500 15960
rect 5776 15920 5782 15932
rect 4709 15895 4767 15901
rect 4709 15861 4721 15895
rect 4755 15861 4767 15895
rect 4709 15855 4767 15861
rect 4798 15852 4804 15904
rect 4856 15892 4862 15904
rect 4893 15895 4951 15901
rect 4893 15892 4905 15895
rect 4856 15864 4905 15892
rect 4856 15852 4862 15864
rect 4893 15861 4905 15864
rect 4939 15861 4951 15895
rect 4893 15855 4951 15861
rect 5353 15895 5411 15901
rect 5353 15861 5365 15895
rect 5399 15892 5411 15895
rect 6362 15892 6368 15904
rect 5399 15864 6368 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6472 15892 6500 15932
rect 8202 15920 8208 15972
rect 8260 15960 8266 15972
rect 8680 15960 8708 16000
rect 9125 15997 9137 16000
rect 9171 15997 9183 16031
rect 9306 16028 9312 16040
rect 9267 16000 9312 16028
rect 9125 15991 9183 15997
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 9398 15988 9404 16040
rect 9456 15988 9462 16040
rect 9674 15988 9680 16040
rect 9732 15988 9738 16040
rect 10152 16037 10180 16068
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 11020 16000 11161 16028
rect 11020 15988 11026 16000
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 8260 15932 8708 15960
rect 9325 15960 9353 15988
rect 10980 15960 11008 15988
rect 9325 15932 11008 15960
rect 8260 15920 8266 15932
rect 8662 15892 8668 15904
rect 6472 15864 8668 15892
rect 8662 15852 8668 15864
rect 8720 15852 8726 15904
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 9398 15892 9404 15904
rect 9180 15864 9404 15892
rect 9180 15852 9186 15864
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 9769 15895 9827 15901
rect 9769 15892 9781 15895
rect 9732 15864 9781 15892
rect 9732 15852 9738 15864
rect 9769 15861 9781 15864
rect 9815 15861 9827 15895
rect 9769 15855 9827 15861
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10597 15895 10655 15901
rect 10597 15892 10609 15895
rect 10468 15864 10609 15892
rect 10468 15852 10474 15864
rect 10597 15861 10609 15864
rect 10643 15861 10655 15895
rect 11256 15892 11284 16068
rect 11348 16037 11376 16136
rect 11333 16031 11391 16037
rect 11333 15997 11345 16031
rect 11379 15997 11391 16031
rect 11333 15991 11391 15997
rect 11606 15988 11612 16040
rect 11664 15988 11670 16040
rect 11716 16037 11744 16204
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 11885 16167 11943 16173
rect 11885 16133 11897 16167
rect 11931 16133 11943 16167
rect 11885 16127 11943 16133
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 16028 11759 16031
rect 11790 16028 11796 16040
rect 11747 16000 11796 16028
rect 11747 15997 11759 16000
rect 11701 15991 11759 15997
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 11514 15920 11520 15972
rect 11572 15920 11578 15972
rect 11900 15960 11928 16127
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12066 16028 12072 16040
rect 12023 16000 12072 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12066 15988 12072 16000
rect 12124 15988 12130 16040
rect 13538 15988 13544 16040
rect 13596 15988 13602 16040
rect 13725 16031 13783 16037
rect 13725 15997 13737 16031
rect 13771 15997 13783 16031
rect 13725 15991 13783 15997
rect 12222 15963 12280 15969
rect 12222 15960 12234 15963
rect 11900 15932 12234 15960
rect 12222 15929 12234 15932
rect 12268 15929 12280 15963
rect 12222 15923 12280 15929
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 13740 15960 13768 15991
rect 12584 15932 13768 15960
rect 12584 15920 12590 15932
rect 13078 15892 13084 15904
rect 11256 15864 13084 15892
rect 10597 15855 10655 15861
rect 13078 15852 13084 15864
rect 13136 15892 13142 15904
rect 13357 15895 13415 15901
rect 13357 15892 13369 15895
rect 13136 15864 13369 15892
rect 13136 15852 13142 15864
rect 13357 15861 13369 15864
rect 13403 15861 13415 15895
rect 13357 15855 13415 15861
rect 13538 15852 13544 15904
rect 13596 15852 13602 15904
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 5902 15648 5908 15700
rect 5960 15688 5966 15700
rect 8478 15688 8484 15700
rect 5960 15660 8484 15688
rect 5960 15648 5966 15660
rect 4982 15580 4988 15632
rect 5040 15620 5046 15632
rect 5813 15623 5871 15629
rect 5813 15620 5825 15623
rect 5040 15592 5825 15620
rect 5040 15580 5046 15592
rect 5813 15589 5825 15592
rect 5859 15589 5871 15623
rect 5813 15583 5871 15589
rect 5994 15580 6000 15632
rect 6052 15580 6058 15632
rect 7668 15629 7696 15660
rect 8478 15648 8484 15660
rect 8536 15688 8542 15700
rect 10226 15688 10232 15700
rect 8536 15660 10232 15688
rect 8536 15648 8542 15660
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 10505 15691 10563 15697
rect 10505 15657 10517 15691
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 7653 15623 7711 15629
rect 7653 15589 7665 15623
rect 7699 15589 7711 15623
rect 7653 15583 7711 15589
rect 7745 15623 7803 15629
rect 7745 15589 7757 15623
rect 7791 15620 7803 15623
rect 8021 15623 8079 15629
rect 8021 15620 8033 15623
rect 7791 15592 8033 15620
rect 7791 15589 7803 15592
rect 7745 15583 7803 15589
rect 8021 15589 8033 15592
rect 8067 15589 8079 15623
rect 10137 15623 10195 15629
rect 8021 15583 8079 15589
rect 8128 15592 9996 15620
rect 8128 15564 8156 15592
rect 2314 15512 2320 15564
rect 2372 15512 2378 15564
rect 2584 15555 2642 15561
rect 2584 15521 2596 15555
rect 2630 15552 2642 15555
rect 3326 15552 3332 15564
rect 2630 15524 3332 15552
rect 2630 15521 2642 15524
rect 2584 15515 2642 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4157 15555 4215 15561
rect 4157 15521 4169 15555
rect 4203 15552 4215 15555
rect 4338 15552 4344 15564
rect 4203 15524 4344 15552
rect 4203 15521 4215 15524
rect 4157 15515 4215 15521
rect 4338 15512 4344 15524
rect 4396 15512 4402 15564
rect 7561 15555 7619 15561
rect 7561 15521 7573 15555
rect 7607 15521 7619 15555
rect 7561 15515 7619 15521
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 8110 15552 8116 15564
rect 7975 15524 8116 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 4246 15444 4252 15496
rect 4304 15444 4310 15496
rect 7576 15484 7604 15515
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9030 15512 9036 15564
rect 9088 15512 9094 15564
rect 9122 15512 9128 15564
rect 9180 15512 9186 15564
rect 9306 15512 9312 15564
rect 9364 15512 9370 15564
rect 9582 15561 9588 15564
rect 9401 15555 9459 15561
rect 9401 15521 9413 15555
rect 9447 15521 9459 15555
rect 9401 15515 9459 15521
rect 9539 15555 9588 15561
rect 9539 15521 9551 15555
rect 9585 15521 9588 15555
rect 9539 15515 9588 15521
rect 7576 15456 7696 15484
rect 3418 15376 3424 15428
rect 3476 15416 3482 15428
rect 3789 15419 3847 15425
rect 3789 15416 3801 15419
rect 3476 15388 3801 15416
rect 3476 15376 3482 15388
rect 3789 15385 3801 15388
rect 3835 15385 3847 15419
rect 7668 15416 7696 15456
rect 8570 15444 8576 15496
rect 8628 15444 8634 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 9141 15484 9169 15512
rect 8720 15456 9169 15484
rect 8720 15444 8726 15456
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 9416 15484 9444 15515
rect 9582 15512 9588 15515
rect 9640 15512 9646 15564
rect 9968 15561 9996 15592
rect 10137 15589 10149 15623
rect 10183 15620 10195 15623
rect 10410 15620 10416 15632
rect 10183 15592 10416 15620
rect 10183 15589 10195 15592
rect 10137 15583 10195 15589
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 10520 15620 10548 15651
rect 10962 15648 10968 15700
rect 11020 15648 11026 15700
rect 11514 15648 11520 15700
rect 11572 15688 11578 15700
rect 12437 15691 12495 15697
rect 12437 15688 12449 15691
rect 11572 15660 12449 15688
rect 11572 15648 11578 15660
rect 12437 15657 12449 15660
rect 12483 15657 12495 15691
rect 12437 15651 12495 15657
rect 12078 15623 12136 15629
rect 12078 15620 12090 15623
rect 10520 15592 12090 15620
rect 12078 15589 12090 15592
rect 12124 15589 12136 15623
rect 12078 15583 12136 15589
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 10226 15512 10232 15564
rect 10284 15512 10290 15564
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15552 10379 15555
rect 10502 15552 10508 15564
rect 10367 15524 10508 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 10502 15512 10508 15524
rect 10560 15552 10566 15564
rect 11238 15552 11244 15564
rect 10560 15524 11244 15552
rect 10560 15512 10566 15524
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 13078 15512 13084 15564
rect 13136 15512 13142 15564
rect 9272 15456 9444 15484
rect 12345 15487 12403 15493
rect 9272 15444 9278 15456
rect 12345 15453 12357 15487
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 8018 15416 8024 15428
rect 7668 15388 8024 15416
rect 3789 15379 3847 15385
rect 8018 15376 8024 15388
rect 8076 15416 8082 15428
rect 11330 15416 11336 15428
rect 8076 15388 11336 15416
rect 8076 15376 8082 15388
rect 11330 15376 11336 15388
rect 11388 15376 11394 15428
rect 3697 15351 3755 15357
rect 3697 15317 3709 15351
rect 3743 15348 3755 15351
rect 4338 15348 4344 15360
rect 3743 15320 4344 15348
rect 3743 15317 3755 15320
rect 3697 15311 3755 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 6181 15351 6239 15357
rect 6181 15348 6193 15351
rect 6052 15320 6193 15348
rect 6052 15308 6058 15320
rect 6181 15317 6193 15320
rect 6227 15317 6239 15351
rect 6181 15311 6239 15317
rect 7374 15308 7380 15360
rect 7432 15308 7438 15360
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12360 15348 12388 15447
rect 12124 15320 12388 15348
rect 12124 15308 12130 15320
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3326 15144 3332 15156
rect 2915 15116 3332 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3326 15104 3332 15116
rect 3384 15104 3390 15156
rect 6086 15104 6092 15156
rect 6144 15144 6150 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 6144 15116 6377 15144
rect 6144 15104 6150 15116
rect 6365 15113 6377 15116
rect 6411 15144 6423 15147
rect 6638 15144 6644 15156
rect 6411 15116 6644 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 6638 15104 6644 15116
rect 6696 15144 6702 15156
rect 6696 15116 8708 15144
rect 6696 15104 6702 15116
rect 6270 14968 6276 15020
rect 6328 15008 6334 15020
rect 6730 15008 6736 15020
rect 6328 14980 6736 15008
rect 6328 14968 6334 14980
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3237 14943 3295 14949
rect 3237 14940 3249 14943
rect 3099 14912 3249 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3237 14909 3249 14912
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3418 14900 3424 14952
rect 3476 14900 3482 14952
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14940 3663 14943
rect 4614 14940 4620 14952
rect 3651 14912 4620 14940
rect 3651 14909 3663 14912
rect 3605 14903 3663 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 4706 14900 4712 14952
rect 4764 14900 4770 14952
rect 4985 14943 5043 14949
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 6288 14940 6316 14968
rect 5031 14912 6316 14940
rect 7000 14943 7058 14949
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 7000 14909 7012 14943
rect 7046 14940 7058 14943
rect 7374 14940 7380 14952
rect 7046 14912 7380 14940
rect 7046 14909 7058 14912
rect 7000 14903 7058 14909
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 8570 14940 8576 14952
rect 8036 14912 8576 14940
rect 5230 14875 5288 14881
rect 5230 14872 5242 14875
rect 4908 14844 5242 14872
rect 4908 14813 4936 14844
rect 5230 14841 5242 14844
rect 5276 14841 5288 14875
rect 5230 14835 5288 14841
rect 4893 14807 4951 14813
rect 4893 14773 4905 14807
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 8036 14804 8064 14912
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 8389 14875 8447 14881
rect 8389 14841 8401 14875
rect 8435 14872 8447 14875
rect 8680 14872 8708 15116
rect 12526 15008 12532 15020
rect 11440 14980 12020 15008
rect 11238 14900 11244 14952
rect 11296 14900 11302 14952
rect 11440 14949 11468 14980
rect 11425 14943 11483 14949
rect 11425 14909 11437 14943
rect 11471 14909 11483 14943
rect 11425 14903 11483 14909
rect 11790 14900 11796 14952
rect 11848 14900 11854 14952
rect 11992 14949 12020 14980
rect 12406 14980 12532 15008
rect 11977 14943 12035 14949
rect 11977 14909 11989 14943
rect 12023 14940 12035 14943
rect 12406 14940 12434 14980
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 12023 14912 12434 14940
rect 12023 14909 12035 14912
rect 11977 14903 12035 14909
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13136 14912 13737 14940
rect 13136 14900 13142 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 13814 14900 13820 14952
rect 13872 14940 13878 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13872 14912 13921 14940
rect 13872 14900 13878 14912
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 8435 14844 8708 14872
rect 8435 14841 8447 14844
rect 8389 14835 8447 14841
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 11885 14875 11943 14881
rect 11885 14872 11897 14875
rect 11204 14844 11897 14872
rect 11204 14832 11210 14844
rect 11885 14841 11897 14844
rect 11931 14841 11943 14875
rect 11885 14835 11943 14841
rect 8113 14807 8171 14813
rect 8113 14804 8125 14807
rect 7432 14776 8125 14804
rect 7432 14764 7438 14776
rect 8113 14773 8125 14776
rect 8159 14773 8171 14807
rect 8113 14767 8171 14773
rect 8202 14764 8208 14816
rect 8260 14804 8266 14816
rect 8757 14807 8815 14813
rect 8757 14804 8769 14807
rect 8260 14776 8769 14804
rect 8260 14764 8266 14776
rect 8757 14773 8769 14776
rect 8803 14773 8815 14807
rect 8757 14767 8815 14773
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 10226 14804 10232 14816
rect 9824 14776 10232 14804
rect 9824 14764 9830 14776
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11698 14804 11704 14816
rect 11379 14776 11704 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11698 14764 11704 14776
rect 11756 14764 11762 14816
rect 13817 14807 13875 14813
rect 13817 14773 13829 14807
rect 13863 14804 13875 14807
rect 13906 14804 13912 14816
rect 13863 14776 13912 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 13906 14764 13912 14776
rect 13964 14764 13970 14816
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 3237 14603 3295 14609
rect 3237 14569 3249 14603
rect 3283 14600 3295 14603
rect 3283 14572 3556 14600
rect 3283 14569 3295 14572
rect 3237 14563 3295 14569
rect 2314 14532 2320 14544
rect 1872 14504 2320 14532
rect 1872 14473 1900 14504
rect 2314 14492 2320 14504
rect 2372 14492 2378 14544
rect 3418 14492 3424 14544
rect 3476 14532 3482 14544
rect 3528 14541 3556 14572
rect 3602 14560 3608 14612
rect 3660 14600 3666 14612
rect 3957 14603 4015 14609
rect 3957 14600 3969 14603
rect 3660 14572 3969 14600
rect 3660 14560 3666 14572
rect 3957 14569 3969 14572
rect 4003 14600 4015 14603
rect 4246 14600 4252 14612
rect 4003 14572 4252 14600
rect 4003 14569 4015 14572
rect 3957 14563 4015 14569
rect 4246 14560 4252 14572
rect 4304 14560 4310 14612
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 4764 14572 5825 14600
rect 4764 14560 4770 14572
rect 5813 14569 5825 14572
rect 5859 14569 5871 14603
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 5813 14563 5871 14569
rect 5920 14572 7021 14600
rect 3513 14535 3571 14541
rect 3513 14532 3525 14535
rect 3476 14504 3525 14532
rect 3476 14492 3482 14504
rect 3513 14501 3525 14504
rect 3559 14501 3571 14535
rect 3513 14495 3571 14501
rect 4157 14535 4215 14541
rect 4157 14501 4169 14535
rect 4203 14532 4215 14535
rect 4614 14532 4620 14544
rect 4203 14504 4620 14532
rect 4203 14501 4215 14504
rect 4157 14495 4215 14501
rect 4614 14492 4620 14504
rect 4672 14532 4678 14544
rect 5920 14532 5948 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7009 14563 7067 14569
rect 11054 14560 11060 14612
rect 11112 14560 11118 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 13630 14600 13636 14612
rect 13495 14572 13636 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 4672 14504 5948 14532
rect 5997 14535 6055 14541
rect 4672 14492 4678 14504
rect 5997 14501 6009 14535
rect 6043 14532 6055 14535
rect 7653 14535 7711 14541
rect 6043 14504 6500 14532
rect 6043 14501 6055 14504
rect 5997 14495 6055 14501
rect 6472 14476 6500 14504
rect 7653 14501 7665 14535
rect 7699 14532 7711 14535
rect 8202 14532 8208 14544
rect 7699 14504 8208 14532
rect 7699 14501 7711 14504
rect 7653 14495 7711 14501
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 8297 14535 8355 14541
rect 8297 14501 8309 14535
rect 8343 14532 8355 14535
rect 8757 14535 8815 14541
rect 8757 14532 8769 14535
rect 8343 14504 8769 14532
rect 8343 14501 8355 14504
rect 8297 14495 8355 14501
rect 8757 14501 8769 14504
rect 8803 14501 8815 14535
rect 13078 14532 13084 14544
rect 8757 14495 8815 14501
rect 9646 14504 11008 14532
rect 2130 14473 2136 14476
rect 1857 14467 1915 14473
rect 1857 14433 1869 14467
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 2124 14427 2136 14473
rect 2130 14424 2136 14427
rect 2188 14424 2194 14476
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 3329 14467 3387 14473
rect 3329 14464 3341 14467
rect 3292 14436 3341 14464
rect 3292 14424 3298 14436
rect 3329 14433 3341 14436
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6362 14464 6368 14476
rect 5960 14436 6368 14464
rect 5960 14424 5966 14436
rect 6362 14424 6368 14436
rect 6420 14424 6426 14476
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 7926 14473 7932 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6512 14436 6929 14464
rect 6512 14424 6518 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 6917 14427 6975 14433
rect 7024 14436 7389 14464
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 7024 14396 7052 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 7470 14467 7528 14473
rect 7470 14433 7482 14467
rect 7516 14433 7528 14467
rect 7470 14427 7528 14433
rect 7745 14467 7803 14473
rect 7745 14433 7757 14467
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 7883 14467 7932 14473
rect 7883 14433 7895 14467
rect 7929 14433 7932 14467
rect 7883 14427 7932 14433
rect 4488 14368 7052 14396
rect 4488 14356 4494 14368
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7484 14396 7512 14427
rect 7340 14368 7512 14396
rect 7760 14396 7788 14427
rect 7926 14424 7932 14427
rect 7984 14424 7990 14476
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 8386 14424 8392 14476
rect 8444 14424 8450 14476
rect 8478 14424 8484 14476
rect 8536 14464 8542 14476
rect 9646 14464 9674 14504
rect 8536 14436 9674 14464
rect 9953 14467 10011 14473
rect 8536 14424 8542 14436
rect 9953 14433 9965 14467
rect 9999 14433 10011 14467
rect 9953 14427 10011 14433
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10318 14464 10324 14476
rect 10183 14436 10324 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 8018 14396 8024 14408
rect 7760 14368 8024 14396
rect 7340 14356 7346 14368
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8404 14396 8432 14424
rect 8404 14368 9352 14396
rect 3697 14331 3755 14337
rect 3697 14297 3709 14331
rect 3743 14328 3755 14331
rect 8665 14331 8723 14337
rect 3743 14300 4016 14328
rect 3743 14297 3755 14300
rect 3697 14291 3755 14297
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 3988 14269 4016 14300
rect 8665 14297 8677 14331
rect 8711 14328 8723 14331
rect 8938 14328 8944 14340
rect 8711 14300 8944 14328
rect 8711 14297 8723 14300
rect 8665 14291 8723 14297
rect 8938 14288 8944 14300
rect 8996 14288 9002 14340
rect 9324 14328 9352 14368
rect 9398 14356 9404 14408
rect 9456 14356 9462 14408
rect 9968 14396 9996 14427
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 10980 14473 11008 14504
rect 11256 14504 13084 14532
rect 11256 14476 11284 14504
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 11238 14424 11244 14476
rect 11296 14424 11302 14476
rect 11330 14424 11336 14476
rect 11388 14464 11394 14476
rect 11425 14467 11483 14473
rect 11425 14464 11437 14467
rect 11388 14436 11437 14464
rect 11388 14424 11394 14436
rect 11425 14433 11437 14436
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 11609 14467 11667 14473
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 12526 14464 12532 14476
rect 11655 14436 12532 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 11624 14396 11652 14427
rect 12526 14424 12532 14436
rect 12584 14464 12590 14476
rect 13354 14464 13360 14476
rect 12584 14436 13360 14464
rect 12584 14424 12590 14436
rect 13354 14424 13360 14436
rect 13412 14424 13418 14476
rect 13906 14473 13912 14476
rect 13900 14464 13912 14473
rect 13867 14436 13912 14464
rect 13900 14427 13912 14436
rect 13906 14424 13912 14427
rect 13964 14424 13970 14476
rect 9968 14368 11652 14396
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 13633 14399 13691 14405
rect 13633 14396 13645 14399
rect 12124 14368 13645 14396
rect 12124 14356 12130 14368
rect 13633 14365 13645 14368
rect 13679 14365 13691 14399
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 13633 14359 13691 14365
rect 15028 14368 15669 14396
rect 9324 14300 12434 14328
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 5994 14220 6000 14272
rect 6052 14220 6058 14272
rect 8021 14263 8079 14269
rect 8021 14229 8033 14263
rect 8067 14260 8079 14263
rect 9214 14260 9220 14272
rect 8067 14232 9220 14260
rect 8067 14229 8079 14232
rect 8021 14223 8079 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 10045 14263 10103 14269
rect 10045 14229 10057 14263
rect 10091 14260 10103 14263
rect 10778 14260 10784 14272
rect 10091 14232 10784 14260
rect 10091 14229 10103 14232
rect 10045 14223 10103 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 12406 14260 12434 14300
rect 14918 14288 14924 14340
rect 14976 14328 14982 14340
rect 15028 14337 15056 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15013 14331 15071 14337
rect 15013 14328 15025 14331
rect 14976 14300 15025 14328
rect 14976 14288 14982 14300
rect 15013 14297 15025 14300
rect 15059 14297 15071 14331
rect 15013 14291 15071 14297
rect 13906 14260 13912 14272
rect 12406 14232 13912 14260
rect 13906 14220 13912 14232
rect 13964 14220 13970 14272
rect 13998 14220 14004 14272
rect 14056 14260 14062 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14056 14232 15117 14260
rect 14056 14220 14062 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 2317 14059 2375 14065
rect 2317 14056 2329 14059
rect 2188 14028 2329 14056
rect 2188 14016 2194 14028
rect 2317 14025 2329 14028
rect 2363 14025 2375 14059
rect 2317 14019 2375 14025
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4019 14028 4200 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 3602 13988 3608 14000
rect 3375 13960 3608 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 3602 13948 3608 13960
rect 3660 13948 3666 14000
rect 4172 13988 4200 14028
rect 4430 14016 4436 14068
rect 4488 14016 4494 14068
rect 5169 14059 5227 14065
rect 5169 14025 5181 14059
rect 5215 14025 5227 14059
rect 5169 14019 5227 14025
rect 5184 13988 5212 14019
rect 7282 14016 7288 14068
rect 7340 14016 7346 14068
rect 7926 14016 7932 14068
rect 7984 14016 7990 14068
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8113 14059 8171 14065
rect 8113 14056 8125 14059
rect 8076 14028 8125 14056
rect 8076 14016 8082 14028
rect 8113 14025 8125 14028
rect 8159 14025 8171 14059
rect 9398 14056 9404 14068
rect 8113 14019 8171 14025
rect 8220 14028 9404 14056
rect 5442 13988 5448 14000
rect 4172 13960 5448 13988
rect 5442 13948 5448 13960
rect 5500 13948 5506 14000
rect 3786 13920 3792 13932
rect 2516 13892 3792 13920
rect 2516 13861 2544 13892
rect 3786 13880 3792 13892
rect 3844 13880 3850 13932
rect 4065 13923 4123 13929
rect 4065 13889 4077 13923
rect 4111 13920 4123 13923
rect 4338 13920 4344 13932
rect 4111 13892 4344 13920
rect 4111 13889 4123 13892
rect 4065 13883 4123 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 8220 13920 8248 14028
rect 9398 14016 9404 14028
rect 9456 14056 9462 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9456 14028 10057 14056
rect 9456 14016 9462 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13814 14056 13820 14068
rect 13587 14028 13820 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 8481 13991 8539 13997
rect 8481 13957 8493 13991
rect 8527 13988 8539 13991
rect 8662 13988 8668 14000
rect 8527 13960 8668 13988
rect 8527 13957 8539 13960
rect 8481 13951 8539 13957
rect 8662 13948 8668 13960
rect 8720 13948 8726 14000
rect 11330 13948 11336 14000
rect 11388 13948 11394 14000
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 11480 13960 12296 13988
rect 11480 13948 11486 13960
rect 12066 13920 12072 13932
rect 7760 13892 8248 13920
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13821 2559 13855
rect 2501 13815 2559 13821
rect 3234 13812 3240 13864
rect 3292 13812 3298 13864
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 3973 13855 4031 13861
rect 3973 13852 3985 13855
rect 3476 13824 3985 13852
rect 3476 13812 3482 13824
rect 3973 13821 3985 13824
rect 4019 13821 4031 13855
rect 3973 13815 4031 13821
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 4212 13824 4261 13852
rect 4212 13812 4218 13824
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 6178 13852 6184 13864
rect 4249 13815 4307 13821
rect 5123 13821 5181 13827
rect 5123 13787 5135 13821
rect 5169 13818 5181 13821
rect 5276 13824 6184 13852
rect 5276 13818 5304 13824
rect 5169 13790 5304 13818
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 6696 13824 7205 13852
rect 6696 13812 6702 13824
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7374 13812 7380 13864
rect 7432 13812 7438 13864
rect 7760 13861 7788 13892
rect 8220 13861 8248 13892
rect 11532 13892 12072 13920
rect 7561 13855 7619 13861
rect 7561 13821 7573 13855
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8021 13855 8079 13861
rect 8021 13821 8033 13855
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 8205 13855 8263 13861
rect 8205 13821 8217 13855
rect 8251 13821 8263 13855
rect 8205 13815 8263 13821
rect 5169 13787 5181 13790
rect 5123 13781 5181 13787
rect 5353 13787 5411 13793
rect 5353 13753 5365 13787
rect 5399 13784 5411 13787
rect 5534 13784 5540 13796
rect 5399 13756 5540 13784
rect 5399 13753 5411 13756
rect 5353 13747 5411 13753
rect 5534 13744 5540 13756
rect 5592 13744 5598 13796
rect 5902 13744 5908 13796
rect 5960 13744 5966 13796
rect 6089 13787 6147 13793
rect 6089 13753 6101 13787
rect 6135 13784 6147 13787
rect 7098 13784 7104 13796
rect 6135 13756 7104 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 7576 13784 7604 13815
rect 8036 13784 8064 13815
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 8352 13824 8401 13852
rect 8352 13812 8358 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8478 13812 8484 13864
rect 8536 13852 8542 13864
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8536 13824 8677 13852
rect 8536 13812 8542 13824
rect 8665 13821 8677 13824
rect 8711 13852 8723 13855
rect 11532 13852 11560 13892
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 12268 13929 12296 13960
rect 13630 13948 13636 14000
rect 13688 13988 13694 14000
rect 13688 13960 14688 13988
rect 13688 13948 13694 13960
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13889 12311 13923
rect 12253 13883 12311 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12952 13892 13093 13920
rect 12952 13880 12958 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13504 13892 13829 13920
rect 13504 13880 13510 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 13998 13920 14004 13932
rect 13817 13883 13875 13889
rect 13924 13892 14004 13920
rect 8711 13824 11560 13852
rect 11609 13855 11667 13861
rect 8711 13821 8723 13824
rect 8665 13815 8723 13821
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 12161 13855 12219 13861
rect 11655 13824 11744 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 8938 13793 8944 13796
rect 8932 13784 8944 13793
rect 7576 13756 8064 13784
rect 8899 13756 8944 13784
rect 4982 13676 4988 13728
rect 5040 13676 5046 13728
rect 6273 13719 6331 13725
rect 6273 13685 6285 13719
rect 6319 13716 6331 13719
rect 6546 13716 6552 13728
rect 6319 13688 6552 13716
rect 6319 13685 6331 13688
rect 6273 13679 6331 13685
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7576 13716 7604 13756
rect 8932 13747 8944 13756
rect 8938 13744 8944 13747
rect 8996 13744 9002 13796
rect 11238 13744 11244 13796
rect 11296 13784 11302 13796
rect 11333 13787 11391 13793
rect 11333 13784 11345 13787
rect 11296 13756 11345 13784
rect 11296 13744 11302 13756
rect 11333 13753 11345 13756
rect 11379 13753 11391 13787
rect 11333 13747 11391 13753
rect 11514 13744 11520 13796
rect 11572 13744 11578 13796
rect 11716 13725 11744 13824
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12802 13852 12808 13864
rect 12207 13824 12808 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13354 13812 13360 13864
rect 13412 13852 13418 13864
rect 13924 13861 13952 13892
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 14660 13861 14688 13960
rect 13909 13855 13967 13861
rect 13412 13824 13860 13852
rect 13412 13812 13418 13824
rect 12069 13787 12127 13793
rect 12069 13753 12081 13787
rect 12115 13784 12127 13787
rect 13832 13784 13860 13824
rect 13909 13821 13921 13855
rect 13955 13821 13967 13855
rect 14185 13855 14243 13861
rect 14185 13852 14197 13855
rect 13909 13815 13967 13821
rect 14016 13824 14197 13852
rect 14016 13784 14044 13824
rect 14185 13821 14197 13824
rect 14231 13821 14243 13855
rect 14185 13815 14243 13821
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 14645 13855 14703 13861
rect 14415 13824 14596 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 12115 13756 13032 13784
rect 13832 13756 14044 13784
rect 14568 13784 14596 13824
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14918 13852 14924 13864
rect 14645 13815 14703 13821
rect 14752 13824 14924 13852
rect 14752 13784 14780 13824
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 14568 13756 14780 13784
rect 12115 13753 12127 13756
rect 12069 13747 12127 13753
rect 13004 13728 13032 13756
rect 6972 13688 7604 13716
rect 11701 13719 11759 13725
rect 6972 13676 6978 13688
rect 11701 13685 11713 13719
rect 11747 13685 11759 13719
rect 11701 13679 11759 13685
rect 12526 13676 12532 13728
rect 12584 13676 12590 13728
rect 12802 13676 12808 13728
rect 12860 13716 12866 13728
rect 12897 13719 12955 13725
rect 12897 13716 12909 13719
rect 12860 13688 12909 13716
rect 12860 13676 12866 13688
rect 12897 13685 12909 13688
rect 12943 13685 12955 13719
rect 12897 13679 12955 13685
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 13630 13716 13636 13728
rect 13044 13688 13636 13716
rect 13044 13676 13050 13688
rect 13630 13676 13636 13688
rect 13688 13716 13694 13728
rect 15028 13716 15056 13815
rect 13688 13688 15056 13716
rect 13688 13676 13694 13688
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2792 13484 3065 13512
rect 2685 13447 2743 13453
rect 2685 13444 2697 13447
rect 2424 13416 2697 13444
rect 2424 13385 2452 13416
rect 2685 13413 2697 13416
rect 2731 13413 2743 13447
rect 2685 13407 2743 13413
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13345 2467 13379
rect 2409 13339 2467 13345
rect 2593 13379 2651 13385
rect 2593 13345 2605 13379
rect 2639 13376 2651 13379
rect 2792 13376 2820 13484
rect 3053 13481 3065 13484
rect 3099 13512 3111 13515
rect 3234 13512 3240 13524
rect 3099 13484 3240 13512
rect 3099 13481 3111 13484
rect 3053 13475 3111 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4893 13515 4951 13521
rect 4893 13512 4905 13515
rect 4663 13484 4905 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4893 13481 4905 13484
rect 4939 13481 4951 13515
rect 5534 13512 5540 13524
rect 4893 13475 4951 13481
rect 5184 13484 5540 13512
rect 2884 13416 3280 13444
rect 2884 13385 2912 13416
rect 3252 13385 3280 13416
rect 2639 13348 2820 13376
rect 2869 13379 2927 13385
rect 2639 13345 2651 13348
rect 2593 13339 2651 13345
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13345 3019 13379
rect 2961 13339 3019 13345
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 3283 13348 4261 13376
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 4249 13345 4261 13348
rect 4295 13376 4307 13379
rect 4982 13376 4988 13388
rect 4295 13348 4988 13376
rect 4295 13345 4307 13348
rect 4249 13339 4307 13345
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2976 13308 3004 13339
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 5184 13385 5212 13484
rect 5534 13472 5540 13484
rect 5592 13512 5598 13524
rect 6914 13512 6920 13524
rect 5592 13484 6920 13512
rect 5592 13472 5598 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 12066 13472 12072 13524
rect 12124 13512 12130 13524
rect 12253 13515 12311 13521
rect 12253 13512 12265 13515
rect 12124 13484 12265 13512
rect 12124 13472 12130 13484
rect 12253 13481 12265 13484
rect 12299 13481 12311 13515
rect 12253 13475 12311 13481
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 14458 13512 14464 13524
rect 12860 13484 14464 13512
rect 12860 13472 12866 13484
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 6454 13404 6460 13456
rect 6512 13444 6518 13456
rect 6549 13447 6607 13453
rect 6549 13444 6561 13447
rect 6512 13416 6561 13444
rect 6512 13404 6518 13416
rect 6549 13413 6561 13416
rect 6595 13444 6607 13447
rect 6638 13444 6644 13456
rect 6595 13416 6644 13444
rect 6595 13413 6607 13416
rect 6549 13407 6607 13413
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 6730 13404 6736 13456
rect 6788 13444 6794 13456
rect 7285 13447 7343 13453
rect 7285 13444 7297 13447
rect 6788 13416 7297 13444
rect 6788 13404 6794 13416
rect 7285 13413 7297 13416
rect 7331 13413 7343 13447
rect 7285 13407 7343 13413
rect 9033 13447 9091 13453
rect 9033 13413 9045 13447
rect 9079 13444 9091 13447
rect 9858 13444 9864 13456
rect 9079 13416 9864 13444
rect 9079 13413 9091 13416
rect 9033 13407 9091 13413
rect 9858 13404 9864 13416
rect 9916 13444 9922 13456
rect 10965 13447 11023 13453
rect 10965 13444 10977 13447
rect 9916 13416 10977 13444
rect 9916 13404 9922 13416
rect 10965 13413 10977 13416
rect 11011 13413 11023 13447
rect 10965 13407 11023 13413
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 5077 13339 5135 13345
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13345 5227 13379
rect 5169 13339 5227 13345
rect 5353 13379 5411 13385
rect 5353 13345 5365 13379
rect 5399 13376 5411 13379
rect 5442 13376 5448 13388
rect 5399 13348 5448 13376
rect 5399 13345 5411 13348
rect 5353 13339 5411 13345
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 2976 13280 3433 13308
rect 2685 13271 2743 13277
rect 3421 13277 3433 13280
rect 3467 13308 3479 13311
rect 3513 13311 3571 13317
rect 3513 13308 3525 13311
rect 3467 13280 3525 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3513 13277 3525 13280
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 2498 13172 2504 13184
rect 2455 13144 2504 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 2700 13172 2728 13271
rect 4154 13268 4160 13320
rect 4212 13268 4218 13320
rect 5092 13308 5120 13339
rect 5442 13336 5448 13348
rect 5500 13336 5506 13388
rect 6178 13336 6184 13388
rect 6236 13376 6242 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6236 13348 6837 13376
rect 6236 13336 6242 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 5261 13311 5319 13317
rect 5092 13280 5212 13308
rect 4614 13172 4620 13184
rect 2700 13144 4620 13172
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4798 13132 4804 13184
rect 4856 13132 4862 13184
rect 5184 13172 5212 13280
rect 5261 13277 5273 13311
rect 5307 13277 5319 13311
rect 5261 13271 5319 13277
rect 5276 13240 5304 13271
rect 5902 13268 5908 13320
rect 5960 13308 5966 13320
rect 7024 13308 7052 13339
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7193 13379 7251 13385
rect 7193 13376 7205 13379
rect 7156 13348 7205 13376
rect 7156 13336 7162 13348
rect 7193 13345 7205 13348
rect 7239 13376 7251 13379
rect 8202 13376 8208 13388
rect 7239 13348 8208 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 5960 13280 7052 13308
rect 5960 13268 5966 13280
rect 6733 13243 6791 13249
rect 5276 13212 6684 13240
rect 5902 13172 5908 13184
rect 5184 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 6656 13172 6684 13212
rect 6733 13209 6745 13243
rect 6779 13240 6791 13243
rect 7098 13240 7104 13252
rect 6779 13212 7104 13240
rect 6779 13209 6791 13212
rect 6733 13203 6791 13209
rect 7098 13200 7104 13212
rect 7156 13200 7162 13252
rect 7208 13172 7236 13339
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9214 13336 9220 13388
rect 9272 13336 9278 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13345 9643 13379
rect 9585 13339 9643 13345
rect 9600 13240 9628 13339
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10137 13379 10195 13385
rect 10137 13376 10149 13379
rect 10008 13348 10149 13376
rect 10008 13336 10014 13348
rect 10137 13345 10149 13348
rect 10183 13376 10195 13379
rect 12618 13376 12624 13388
rect 10183 13348 12624 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13170 13336 13176 13388
rect 13228 13376 13234 13388
rect 13449 13379 13507 13385
rect 13449 13376 13461 13379
rect 13228 13348 13461 13376
rect 13228 13336 13234 13348
rect 13449 13345 13461 13348
rect 13495 13345 13507 13379
rect 13449 13339 13507 13345
rect 13630 13336 13636 13388
rect 13688 13336 13694 13388
rect 13722 13336 13728 13388
rect 13780 13336 13786 13388
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 13906 13376 13912 13388
rect 13863 13348 13912 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 13906 13336 13912 13348
rect 13964 13336 13970 13388
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 9766 13308 9772 13320
rect 9723 13280 9772 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 9766 13268 9772 13280
rect 9824 13268 9830 13320
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 10042 13308 10048 13320
rect 9907 13280 10048 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10594 13308 10600 13320
rect 10152 13280 10600 13308
rect 10152 13240 10180 13280
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 9600 13212 10180 13240
rect 6656 13144 7236 13172
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 10284 13144 10333 13172
rect 10284 13132 10290 13144
rect 10321 13141 10333 13144
rect 10367 13172 10379 13175
rect 10962 13172 10968 13184
rect 10367 13144 10968 13172
rect 10367 13141 10379 13144
rect 10321 13135 10379 13141
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 16666 13172 16672 13184
rect 14139 13144 16672 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5442 12968 5448 12980
rect 5215 12940 5448 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 8202 12928 8208 12980
rect 8260 12928 8266 12980
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9456 12940 9689 12968
rect 9456 12928 9462 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 10134 12968 10140 12980
rect 9677 12931 9735 12937
rect 9876 12940 10140 12968
rect 9692 12900 9720 12931
rect 9766 12900 9772 12912
rect 9692 12872 9772 12900
rect 9766 12860 9772 12872
rect 9824 12860 9830 12912
rect 2314 12792 2320 12844
rect 2372 12832 2378 12844
rect 3786 12832 3792 12844
rect 2372 12804 3792 12832
rect 2372 12792 2378 12804
rect 3786 12792 3792 12804
rect 3844 12792 3850 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 9876 12841 9904 12940
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 11514 12968 11520 12980
rect 10428 12940 11520 12968
rect 10318 12860 10324 12912
rect 10376 12860 10382 12912
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6788 12804 6837 12832
rect 6788 12792 6794 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 5537 12767 5595 12773
rect 5537 12764 5549 12767
rect 4672 12736 5549 12764
rect 4672 12724 4678 12736
rect 5537 12733 5549 12736
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12764 6055 12767
rect 6178 12764 6184 12776
rect 6043 12736 6184 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 6178 12724 6184 12736
rect 6236 12724 6242 12776
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12764 6699 12767
rect 6914 12764 6920 12776
rect 6687 12736 6920 12764
rect 6687 12733 6699 12736
rect 6641 12727 6699 12733
rect 4056 12699 4114 12705
rect 4056 12665 4068 12699
rect 4102 12696 4114 12699
rect 4246 12696 4252 12708
rect 4102 12668 4252 12696
rect 4102 12665 4114 12668
rect 4056 12659 4114 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 5905 12699 5963 12705
rect 5905 12665 5917 12699
rect 5951 12696 5963 12699
rect 6656 12696 6684 12727
rect 6914 12724 6920 12736
rect 6972 12724 6978 12776
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12764 9643 12767
rect 9631 12760 9904 12764
rect 9950 12760 9956 12776
rect 9631 12736 9956 12760
rect 9631 12733 9643 12736
rect 9585 12727 9643 12733
rect 9876 12732 9956 12736
rect 9950 12724 9956 12732
rect 10008 12724 10014 12776
rect 10042 12724 10048 12776
rect 10100 12764 10106 12776
rect 10100 12736 10145 12764
rect 10100 12724 10106 12736
rect 10226 12724 10232 12776
rect 10284 12764 10290 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10284 12736 10333 12764
rect 10284 12724 10290 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10428 12764 10456 12940
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11606 12928 11612 12980
rect 11664 12968 11670 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 11664 12940 12173 12968
rect 11664 12928 11670 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 10686 12860 10692 12912
rect 10744 12860 10750 12912
rect 11790 12860 11796 12912
rect 11848 12860 11854 12912
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 12342 12900 12348 12912
rect 12032 12872 12348 12900
rect 12032 12860 12038 12872
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 13081 12903 13139 12909
rect 13081 12869 13093 12903
rect 13127 12900 13139 12903
rect 15102 12900 15108 12912
rect 13127 12872 15108 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 12526 12832 12532 12844
rect 12084 12804 12532 12832
rect 12084 12773 12112 12804
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 10689 12767 10747 12773
rect 10428 12742 10548 12764
rect 10581 12745 10639 12751
rect 10581 12742 10593 12745
rect 10428 12736 10593 12742
rect 10321 12727 10379 12733
rect 10520 12714 10593 12736
rect 10581 12711 10593 12714
rect 10627 12711 10639 12745
rect 10689 12733 10701 12767
rect 10735 12766 10747 12767
rect 10873 12767 10931 12773
rect 10735 12738 10824 12766
rect 10735 12733 10747 12738
rect 10689 12727 10747 12733
rect 5951 12668 6684 12696
rect 7092 12699 7150 12705
rect 5951 12665 5963 12668
rect 5905 12659 5963 12665
rect 7092 12665 7104 12699
rect 7138 12696 7150 12699
rect 7282 12696 7288 12708
rect 7138 12668 7288 12696
rect 7138 12665 7150 12668
rect 7092 12659 7150 12665
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 9490 12696 9496 12708
rect 7392 12668 9496 12696
rect 5810 12588 5816 12640
rect 5868 12588 5874 12640
rect 6089 12631 6147 12637
rect 6089 12597 6101 12631
rect 6135 12628 6147 12631
rect 6178 12628 6184 12640
rect 6135 12600 6184 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 7392 12628 7420 12668
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 10581 12705 10639 12711
rect 10796 12640 10824 12738
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 10888 12696 10916 12727
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 12434 12724 12440 12776
rect 12492 12724 12498 12776
rect 13078 12724 13084 12776
rect 13136 12724 13142 12776
rect 13357 12767 13415 12773
rect 13357 12733 13369 12767
rect 13403 12764 13415 12767
rect 13814 12764 13820 12776
rect 13403 12736 13820 12764
rect 13403 12733 13415 12736
rect 13357 12727 13415 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 10962 12696 10968 12708
rect 10888 12668 10968 12696
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 11793 12699 11851 12705
rect 11793 12696 11805 12699
rect 11020 12668 11805 12696
rect 11020 12656 11026 12668
rect 11793 12665 11805 12668
rect 11839 12696 11851 12699
rect 12161 12699 12219 12705
rect 12161 12696 12173 12699
rect 11839 12668 12173 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 12161 12665 12173 12668
rect 12207 12696 12219 12699
rect 13096 12696 13124 12724
rect 12207 12668 13124 12696
rect 13265 12699 13323 12705
rect 12207 12665 12219 12668
rect 12161 12659 12219 12665
rect 13265 12665 13277 12699
rect 13311 12696 13323 12699
rect 13538 12696 13544 12708
rect 13311 12668 13544 12696
rect 13311 12665 13323 12668
rect 13265 12659 13323 12665
rect 13538 12656 13544 12668
rect 13596 12656 13602 12708
rect 6696 12600 7420 12628
rect 10229 12631 10287 12637
rect 6696 12588 6702 12600
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10410 12628 10416 12640
rect 10275 12600 10416 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 10505 12631 10563 12637
rect 10505 12597 10517 12631
rect 10551 12628 10563 12631
rect 10594 12628 10600 12640
rect 10551 12600 10600 12628
rect 10551 12597 10563 12600
rect 10505 12591 10563 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10778 12588 10784 12640
rect 10836 12588 10842 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 11977 12631 12035 12637
rect 11977 12628 11989 12631
rect 11756 12600 11989 12628
rect 11756 12588 11762 12600
rect 11977 12597 11989 12600
rect 12023 12597 12035 12631
rect 11977 12591 12035 12597
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 4154 12424 4160 12436
rect 3651 12396 4160 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4246 12384 4252 12436
rect 4304 12384 4310 12436
rect 6914 12384 6920 12436
rect 6972 12424 6978 12436
rect 7193 12427 7251 12433
rect 7193 12424 7205 12427
rect 6972 12396 7205 12424
rect 6972 12384 6978 12396
rect 7193 12393 7205 12396
rect 7239 12393 7251 12427
rect 7193 12387 7251 12393
rect 7282 12384 7288 12436
rect 7340 12384 7346 12436
rect 10336 12396 11008 12424
rect 10336 12365 10364 12396
rect 10980 12368 11008 12396
rect 11146 12384 11152 12436
rect 11204 12384 11210 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12393 11391 12427
rect 11333 12387 11391 12393
rect 10321 12359 10379 12365
rect 10321 12325 10333 12359
rect 10367 12325 10379 12359
rect 10321 12319 10379 12325
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 10778 12356 10784 12368
rect 10551 12328 10784 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 10962 12316 10968 12368
rect 11020 12316 11026 12368
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2314 12288 2320 12300
rect 2271 12260 2320 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 2498 12297 2504 12300
rect 2492 12288 2504 12297
rect 2459 12260 2504 12288
rect 2492 12251 2504 12260
rect 2498 12248 2504 12251
rect 2556 12248 2562 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12288 4491 12291
rect 4798 12288 4804 12300
rect 4479 12260 4804 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4798 12248 4804 12260
rect 4856 12248 4862 12300
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6069 12291 6127 12297
rect 6069 12288 6081 12291
rect 5776 12260 6081 12288
rect 5776 12248 5782 12260
rect 6069 12257 6081 12260
rect 6115 12257 6127 12291
rect 6069 12251 6127 12257
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7156 12260 7481 12288
rect 7156 12248 7162 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 10594 12248 10600 12300
rect 10652 12248 10658 12300
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 11348 12288 11376 12387
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 12161 12427 12219 12433
rect 12161 12424 12173 12427
rect 11572 12396 12173 12424
rect 11572 12384 11578 12396
rect 12161 12393 12173 12396
rect 12207 12393 12219 12427
rect 12161 12387 12219 12393
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 12492 12396 13001 12424
rect 12492 12384 12498 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 13814 12384 13820 12436
rect 13872 12384 13878 12436
rect 14277 12427 14335 12433
rect 14277 12393 14289 12427
rect 14323 12424 14335 12427
rect 14458 12424 14464 12436
rect 14323 12396 14464 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 11793 12359 11851 12365
rect 11793 12325 11805 12359
rect 11839 12356 11851 12359
rect 12618 12356 12624 12368
rect 11839 12328 12624 12356
rect 11839 12325 11851 12328
rect 11793 12319 11851 12325
rect 12618 12316 12624 12328
rect 12676 12356 12682 12368
rect 13449 12359 13507 12365
rect 13449 12356 13461 12359
rect 12676 12328 13461 12356
rect 12676 12316 12682 12328
rect 13449 12325 13461 12328
rect 13495 12356 13507 12359
rect 14292 12356 14320 12387
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 13495 12328 14320 12356
rect 13495 12325 13507 12328
rect 13449 12319 13507 12325
rect 11287 12260 11376 12288
rect 11701 12291 11759 12297
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 12526 12288 12532 12300
rect 11747 12260 12532 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 12526 12248 12532 12260
rect 12584 12288 12590 12300
rect 12986 12288 12992 12300
rect 12584 12260 12992 12288
rect 12584 12248 12590 12260
rect 12986 12248 12992 12260
rect 13044 12288 13050 12300
rect 13357 12291 13415 12297
rect 13357 12288 13369 12291
rect 13044 12260 13369 12288
rect 13044 12248 13050 12260
rect 13357 12257 13369 12260
rect 13403 12288 13415 12291
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13403 12260 14197 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 5828 12084 5856 12183
rect 11882 12180 11888 12232
rect 11940 12180 11946 12232
rect 12710 12180 12716 12232
rect 12768 12180 12774 12232
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12189 14427 12223
rect 14369 12183 14427 12189
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 13814 12152 13820 12164
rect 6880 12124 13820 12152
rect 6880 12112 6886 12124
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14384 12152 14412 12183
rect 14056 12124 14412 12152
rect 14056 12112 14062 12124
rect 6730 12084 6736 12096
rect 5828 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 10321 12087 10379 12093
rect 10321 12084 10333 12087
rect 10284 12056 10333 12084
rect 10284 12044 10290 12056
rect 10321 12053 10333 12056
rect 10367 12053 10379 12087
rect 10321 12047 10379 12053
rect 10962 12044 10968 12096
rect 11020 12044 11026 12096
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 5718 11840 5724 11892
rect 5776 11840 5782 11892
rect 6086 11840 6092 11892
rect 6144 11840 6150 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11609 11883 11667 11889
rect 11609 11880 11621 11883
rect 10652 11852 11621 11880
rect 10652 11840 10658 11852
rect 11609 11849 11621 11852
rect 11655 11849 11667 11883
rect 11609 11843 11667 11849
rect 13173 11883 13231 11889
rect 13173 11849 13185 11883
rect 13219 11880 13231 11883
rect 13262 11880 13268 11892
rect 13219 11852 13268 11880
rect 13219 11849 13231 11852
rect 13173 11843 13231 11849
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13446 11840 13452 11892
rect 13504 11880 13510 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13504 11852 13553 11880
rect 13504 11840 13510 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 10686 11812 10692 11824
rect 10376 11784 10692 11812
rect 10376 11772 10382 11784
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12124 11784 14412 11812
rect 12124 11772 12130 11784
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6788 11716 6837 11744
rect 6788 11704 6794 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12434 11744 12440 11756
rect 12299 11716 12440 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 14384 11753 14412 11784
rect 14369 11747 14427 11753
rect 12912 11716 13952 11744
rect 5902 11636 5908 11688
rect 5960 11636 5966 11688
rect 6178 11636 6184 11688
rect 6236 11636 6242 11688
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 6288 11648 9321 11676
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 6288 11608 6316 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9490 11636 9496 11688
rect 9548 11636 9554 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10318 11676 10324 11688
rect 9723 11648 10324 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11676 12127 11679
rect 12618 11676 12624 11688
rect 12115 11648 12624 11676
rect 12115 11645 12127 11648
rect 12069 11639 12127 11645
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 5500 11580 6316 11608
rect 5500 11568 5506 11580
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7070 11611 7128 11617
rect 7070 11608 7082 11611
rect 6972 11580 7082 11608
rect 6972 11568 6978 11580
rect 7070 11577 7082 11580
rect 7116 11577 7128 11611
rect 11790 11608 11796 11620
rect 7070 11571 7128 11577
rect 8220 11580 11796 11608
rect 8220 11549 8248 11580
rect 11790 11568 11796 11580
rect 11848 11568 11854 11620
rect 11977 11611 12035 11617
rect 11977 11577 11989 11611
rect 12023 11608 12035 11611
rect 12023 11580 12204 11608
rect 12023 11577 12035 11580
rect 11977 11571 12035 11577
rect 8205 11543 8263 11549
rect 8205 11509 8217 11543
rect 8251 11509 8263 11543
rect 12176 11540 12204 11580
rect 12250 11568 12256 11620
rect 12308 11608 12314 11620
rect 12912 11608 12940 11716
rect 13170 11636 13176 11688
rect 13228 11636 13234 11688
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13924 11685 13952 11716
rect 14369 11713 14381 11747
rect 14415 11713 14427 11747
rect 14369 11707 14427 11713
rect 13909 11679 13967 11685
rect 13320 11648 13860 11676
rect 13320 11636 13326 11648
rect 12308 11580 12940 11608
rect 12989 11611 13047 11617
rect 12308 11568 12314 11580
rect 12989 11577 13001 11611
rect 13035 11608 13047 11611
rect 13188 11608 13216 11636
rect 13446 11608 13452 11620
rect 13035 11580 13216 11608
rect 13280 11580 13452 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 12526 11540 12532 11552
rect 12176 11512 12532 11540
rect 8205 11503 8263 11509
rect 12526 11500 12532 11512
rect 12584 11500 12590 11552
rect 13194 11543 13252 11549
rect 13194 11509 13206 11543
rect 13240 11540 13252 11543
rect 13280 11540 13308 11580
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 13722 11568 13728 11620
rect 13780 11568 13786 11620
rect 13832 11608 13860 11648
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 13955 11648 14013 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14001 11639 14059 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 14274 11676 14280 11688
rect 14231 11648 14280 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 14274 11636 14280 11648
rect 14332 11636 14338 11688
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 13832 11580 14105 11608
rect 14093 11577 14105 11580
rect 14139 11577 14151 11611
rect 14093 11571 14151 11577
rect 14458 11568 14464 11620
rect 14516 11608 14522 11620
rect 14614 11611 14672 11617
rect 14614 11608 14626 11611
rect 14516 11580 14626 11608
rect 14516 11568 14522 11580
rect 14614 11577 14626 11580
rect 14660 11577 14672 11611
rect 14614 11571 14672 11577
rect 13240 11512 13308 11540
rect 13357 11543 13415 11549
rect 13240 11509 13252 11512
rect 13194 11503 13252 11509
rect 13357 11509 13369 11543
rect 13403 11540 13415 11543
rect 14366 11540 14372 11552
rect 13403 11512 14372 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14918 11500 14924 11552
rect 14976 11540 14982 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 14976 11512 15761 11540
rect 14976 11500 14982 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 15749 11503 15807 11509
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 5261 11339 5319 11345
rect 5261 11305 5273 11339
rect 5307 11336 5319 11339
rect 6822 11336 6828 11348
rect 5307 11308 6828 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 10318 11336 10324 11348
rect 10100 11308 10324 11336
rect 10100 11296 10106 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 10689 11339 10747 11345
rect 10689 11305 10701 11339
rect 10735 11336 10747 11339
rect 10870 11336 10876 11348
rect 10735 11308 10876 11336
rect 10735 11305 10747 11308
rect 10689 11299 10747 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 11882 11296 11888 11348
rect 11940 11296 11946 11348
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 13722 11336 13728 11348
rect 12299 11308 13728 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 10413 11271 10471 11277
rect 10183 11237 10241 11243
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3844 11172 3893 11200
rect 3844 11160 3850 11172
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4137 11203 4195 11209
rect 4137 11200 4149 11203
rect 4028 11172 4149 11200
rect 4028 11160 4034 11172
rect 4137 11169 4149 11172
rect 4183 11169 4195 11203
rect 4137 11163 4195 11169
rect 8478 11160 8484 11212
rect 8536 11160 8542 11212
rect 8754 11209 8760 11212
rect 8748 11163 8760 11209
rect 8754 11160 8760 11163
rect 8812 11160 8818 11212
rect 10183 11203 10195 11237
rect 10229 11234 10241 11237
rect 10413 11237 10425 11271
rect 10459 11268 10471 11271
rect 10505 11271 10563 11277
rect 10505 11268 10517 11271
rect 10459 11240 10517 11268
rect 10459 11237 10471 11240
rect 10229 11203 10256 11234
rect 10413 11231 10471 11237
rect 10505 11237 10517 11240
rect 10551 11268 10563 11271
rect 11238 11268 11244 11280
rect 10551 11240 11244 11268
rect 10551 11237 10563 11240
rect 10505 11231 10563 11237
rect 11238 11228 11244 11240
rect 11296 11228 11302 11280
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 11848 11240 12388 11268
rect 11848 11228 11854 11240
rect 10183 11200 10256 11203
rect 10778 11200 10784 11212
rect 10183 11197 10784 11200
rect 10228 11172 10784 11197
rect 10778 11160 10784 11172
rect 10836 11200 10842 11212
rect 11054 11200 11060 11212
rect 10836 11172 11060 11200
rect 10836 11160 10842 11172
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 12066 11160 12072 11212
rect 12124 11160 12130 11212
rect 12360 11209 12388 11240
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 13446 11160 13452 11212
rect 13504 11160 13510 11212
rect 13556 11200 13584 11308
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 13998 11296 14004 11348
rect 14056 11296 14062 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14553 11339 14611 11345
rect 14553 11336 14565 11339
rect 14516 11308 14565 11336
rect 14516 11296 14522 11308
rect 14553 11305 14565 11308
rect 14599 11305 14611 11339
rect 14553 11299 14611 11305
rect 13633 11271 13691 11277
rect 13633 11237 13645 11271
rect 13679 11268 13691 11271
rect 15838 11268 15844 11280
rect 13679 11240 15844 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 13725 11203 13783 11209
rect 13725 11200 13737 11203
rect 13556 11172 13737 11200
rect 13725 11169 13737 11172
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 13740 11132 13768 11163
rect 13814 11160 13820 11212
rect 13872 11160 13878 11212
rect 14366 11160 14372 11212
rect 14424 11160 14430 11212
rect 14274 11132 14280 11144
rect 13740 11104 14280 11132
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 9490 11024 9496 11076
rect 9548 11064 9554 11076
rect 10505 11067 10563 11073
rect 10505 11064 10517 11067
rect 9548 11036 10517 11064
rect 9548 11024 9554 11036
rect 10505 11033 10517 11036
rect 10551 11033 10563 11067
rect 10505 11027 10563 11033
rect 9858 10956 9864 11008
rect 9916 10956 9922 11008
rect 10229 10999 10287 11005
rect 10229 10965 10241 10999
rect 10275 10996 10287 10999
rect 10318 10996 10324 11008
rect 10275 10968 10324 10996
rect 10275 10965 10287 10968
rect 10229 10959 10287 10965
rect 10318 10956 10324 10968
rect 10376 10996 10382 11008
rect 10870 10996 10876 11008
rect 10376 10968 10876 10996
rect 10376 10956 10382 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 12250 10996 12256 11008
rect 11480 10968 12256 10996
rect 11480 10956 11486 10968
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 4028 10764 4077 10792
rect 4028 10752 4034 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 4982 10752 4988 10804
rect 5040 10792 5046 10804
rect 5040 10764 6868 10792
rect 5040 10752 5046 10764
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 5537 10727 5595 10733
rect 5537 10724 5549 10727
rect 3844 10696 5549 10724
rect 3844 10684 3850 10696
rect 5537 10693 5549 10696
rect 5583 10724 5595 10727
rect 6178 10724 6184 10736
rect 5583 10696 6184 10724
rect 5583 10693 5595 10696
rect 5537 10687 5595 10693
rect 6178 10684 6184 10696
rect 6236 10684 6242 10736
rect 6840 10724 6868 10764
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 8754 10752 8760 10804
rect 8812 10792 8818 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8812 10764 8861 10792
rect 8812 10752 8818 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9490 10752 9496 10804
rect 9548 10752 9554 10804
rect 10336 10764 12434 10792
rect 8478 10724 8484 10736
rect 6840 10696 8484 10724
rect 8478 10684 8484 10696
rect 8536 10724 8542 10736
rect 10137 10727 10195 10733
rect 10137 10724 10149 10727
rect 8536 10696 10149 10724
rect 8536 10684 8542 10696
rect 10137 10693 10149 10696
rect 10183 10693 10195 10727
rect 10137 10687 10195 10693
rect 4522 10616 4528 10668
rect 4580 10616 4586 10668
rect 4982 10616 4988 10668
rect 5040 10616 5046 10668
rect 6365 10659 6423 10665
rect 6365 10625 6377 10659
rect 6411 10656 6423 10659
rect 7650 10656 7656 10668
rect 6411 10628 7656 10656
rect 6411 10625 6423 10628
rect 6365 10619 6423 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 10042 10656 10048 10668
rect 9631 10628 10048 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 4028 10560 4261 10588
rect 4028 10548 4034 10560
rect 4249 10557 4261 10560
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10557 4399 10591
rect 4341 10551 4399 10557
rect 4356 10520 4384 10551
rect 4614 10548 4620 10600
rect 4672 10548 4678 10600
rect 5077 10591 5135 10597
rect 5077 10557 5089 10591
rect 5123 10588 5135 10591
rect 5534 10588 5540 10600
rect 5123 10560 5540 10588
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 6273 10591 6331 10597
rect 6273 10557 6285 10591
rect 6319 10588 6331 10591
rect 6638 10588 6644 10600
rect 6319 10560 6644 10588
rect 6319 10557 6331 10560
rect 6273 10551 6331 10557
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 6730 10548 6736 10600
rect 6788 10548 6794 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 7098 10588 7104 10600
rect 7055 10560 7104 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 7466 10548 7472 10600
rect 7524 10548 7530 10600
rect 9309 10591 9367 10597
rect 9309 10557 9321 10591
rect 9355 10588 9367 10591
rect 9398 10588 9404 10600
rect 9355 10560 9404 10588
rect 9355 10557 9367 10560
rect 9309 10551 9367 10557
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 10336 10597 10364 10764
rect 11057 10727 11115 10733
rect 11057 10724 11069 10727
rect 10612 10696 11069 10724
rect 10321 10591 10379 10597
rect 10321 10557 10333 10591
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10410 10548 10416 10600
rect 10468 10548 10474 10600
rect 10612 10597 10640 10696
rect 11057 10693 11069 10696
rect 11103 10693 11115 10727
rect 12406 10724 12434 10764
rect 12406 10696 15516 10724
rect 11057 10687 11115 10693
rect 13170 10656 13176 10668
rect 11072 10628 13176 10656
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 6362 10520 6368 10532
rect 4356 10492 6368 10520
rect 6362 10480 6368 10492
rect 6420 10480 6426 10532
rect 7653 10523 7711 10529
rect 7653 10520 7665 10523
rect 6748 10492 7665 10520
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5169 10455 5227 10461
rect 5169 10452 5181 10455
rect 4856 10424 5181 10452
rect 4856 10412 4862 10424
rect 5169 10421 5181 10424
rect 5215 10452 5227 10455
rect 5442 10452 5448 10464
rect 5215 10424 5448 10452
rect 5215 10421 5227 10424
rect 5169 10415 5227 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6748 10461 6776 10492
rect 7653 10489 7665 10492
rect 7699 10489 7711 10523
rect 7653 10483 7711 10489
rect 8941 10523 8999 10529
rect 8941 10489 8953 10523
rect 8987 10520 8999 10523
rect 9125 10523 9183 10529
rect 9125 10520 9137 10523
rect 8987 10492 9137 10520
rect 8987 10489 8999 10492
rect 8941 10483 8999 10489
rect 9125 10489 9137 10492
rect 9171 10489 9183 10523
rect 9125 10483 9183 10489
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 10704 10520 10732 10551
rect 10778 10548 10784 10600
rect 10836 10548 10842 10600
rect 10870 10548 10876 10600
rect 10928 10548 10934 10600
rect 11072 10597 11100 10628
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 15488 10665 15516 10696
rect 15473 10659 15531 10665
rect 15473 10625 15485 10659
rect 15519 10656 15531 10659
rect 16206 10656 16212 10668
rect 15519 10628 16212 10656
rect 15519 10625 15531 10628
rect 15473 10619 15531 10625
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10557 11207 10591
rect 13188 10588 13216 10616
rect 15010 10588 15016 10600
rect 13188 10560 15016 10588
rect 11149 10551 11207 10557
rect 10560 10492 10732 10520
rect 10560 10480 10566 10492
rect 6733 10455 6791 10461
rect 6733 10421 6745 10455
rect 6779 10421 6791 10455
rect 6733 10415 6791 10421
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 8018 10452 8024 10464
rect 7064 10424 8024 10452
rect 7064 10412 7070 10424
rect 8018 10412 8024 10424
rect 8076 10412 8082 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10962 10452 10968 10464
rect 9916 10424 10968 10452
rect 9916 10412 9922 10424
rect 10962 10412 10968 10424
rect 11020 10452 11026 10464
rect 11164 10452 11192 10551
rect 15010 10548 15016 10560
rect 15068 10588 15074 10600
rect 15378 10588 15384 10600
rect 15068 10560 15384 10588
rect 15068 10548 15074 10560
rect 15378 10548 15384 10560
rect 15436 10588 15442 10600
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 15436 10560 15577 10588
rect 15436 10548 15442 10560
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15565 10551 15623 10557
rect 15948 10560 16037 10588
rect 11020 10424 11192 10452
rect 11020 10412 11026 10424
rect 11238 10412 11244 10464
rect 11296 10452 11302 10464
rect 11882 10452 11888 10464
rect 11296 10424 11888 10452
rect 11296 10412 11302 10424
rect 11882 10412 11888 10424
rect 11940 10412 11946 10464
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 13722 10452 13728 10464
rect 13044 10424 13728 10452
rect 13044 10412 13050 10424
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 15948 10461 15976 10560
rect 16025 10557 16037 10560
rect 16071 10557 16083 10591
rect 16025 10551 16083 10557
rect 15933 10455 15991 10461
rect 15933 10421 15945 10455
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16022 10412 16028 10464
rect 16080 10452 16086 10464
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 16080 10424 16129 10452
rect 16080 10412 16086 10424
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16117 10415 16175 10421
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 3786 10208 3792 10260
rect 3844 10257 3850 10260
rect 3844 10251 3863 10257
rect 3851 10217 3863 10251
rect 3844 10211 3863 10217
rect 3844 10208 3850 10211
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 4028 10220 4384 10248
rect 4028 10208 4034 10220
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10149 3663 10183
rect 4356 10180 4384 10220
rect 5000 10220 5580 10248
rect 4356 10152 4752 10180
rect 3605 10143 3663 10149
rect 3620 10044 3648 10143
rect 4246 10072 4252 10124
rect 4304 10072 4310 10124
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 4430 10072 4436 10124
rect 4488 10112 4494 10124
rect 4525 10115 4583 10121
rect 4525 10112 4537 10115
rect 4488 10084 4537 10112
rect 4488 10072 4494 10084
rect 4525 10081 4537 10084
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4617 10115 4675 10121
rect 4617 10081 4629 10115
rect 4663 10110 4675 10115
rect 4724 10110 4752 10152
rect 4663 10082 4752 10110
rect 4663 10081 4675 10082
rect 4617 10075 4675 10081
rect 5000 10053 5028 10220
rect 5552 10180 5580 10220
rect 6730 10208 6736 10260
rect 6788 10208 6794 10260
rect 7374 10248 7380 10260
rect 7116 10220 7380 10248
rect 5552 10152 6408 10180
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 3620 10016 4997 10044
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 5276 10044 5304 10075
rect 5350 10072 5356 10124
rect 5408 10072 5414 10124
rect 5552 10121 5580 10152
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10081 6331 10115
rect 6380 10112 6408 10152
rect 7116 10121 7144 10220
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7466 10208 7472 10260
rect 7524 10208 7530 10260
rect 7650 10208 7656 10260
rect 7708 10208 7714 10260
rect 8294 10248 8300 10260
rect 7760 10220 8300 10248
rect 7760 10180 7788 10220
rect 8294 10208 8300 10220
rect 8352 10208 8358 10260
rect 11977 10251 12035 10257
rect 11977 10217 11989 10251
rect 12023 10248 12035 10251
rect 12066 10248 12072 10260
rect 12023 10220 12072 10248
rect 12023 10217 12035 10220
rect 11977 10211 12035 10217
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 13504 10220 13645 10248
rect 13504 10208 13510 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 13740 10220 15332 10248
rect 8386 10180 8392 10192
rect 7208 10152 7788 10180
rect 7852 10152 8392 10180
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6380 10084 6561 10112
rect 6273 10075 6331 10081
rect 6549 10081 6561 10084
rect 6595 10112 6607 10115
rect 7101 10115 7159 10121
rect 7101 10112 7113 10115
rect 6595 10084 7113 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 7101 10081 7113 10084
rect 7147 10081 7159 10115
rect 7101 10075 7159 10081
rect 6178 10044 6184 10056
rect 5276 10016 6184 10044
rect 4985 10007 5043 10013
rect 6178 10004 6184 10016
rect 6236 10044 6242 10056
rect 6288 10044 6316 10075
rect 6236 10016 6316 10044
rect 6457 10047 6515 10053
rect 6236 10004 6242 10016
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 4430 9936 4436 9988
rect 4488 9976 4494 9988
rect 5074 9976 5080 9988
rect 4488 9948 5080 9976
rect 4488 9936 4494 9948
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5442 9936 5448 9988
rect 5500 9936 5506 9988
rect 5534 9936 5540 9988
rect 5592 9976 5598 9988
rect 6472 9976 6500 10007
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 7208 10053 7236 10152
rect 7852 10121 7880 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 12710 10180 12716 10192
rect 12268 10152 12716 10180
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10081 7987 10115
rect 7929 10075 7987 10081
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10013 7251 10047
rect 7193 10007 7251 10013
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7944 10044 7972 10075
rect 8110 10072 8116 10124
rect 8168 10072 8174 10124
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8260 10084 9137 10112
rect 8260 10072 8266 10084
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 8754 10044 8760 10056
rect 7331 10016 8760 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 5592 9948 6500 9976
rect 5592 9936 5598 9948
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4065 9911 4123 9917
rect 4065 9908 4077 9911
rect 3936 9880 4077 9908
rect 3936 9868 3942 9880
rect 4065 9877 4077 9880
rect 4111 9877 4123 9911
rect 4065 9871 4123 9877
rect 4706 9868 4712 9920
rect 4764 9868 4770 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5552 9908 5580 9936
rect 5215 9880 5580 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 6472 9908 6500 9948
rect 6822 9908 6828 9920
rect 6472 9880 6828 9908
rect 6822 9868 6828 9880
rect 6880 9908 6886 9920
rect 7300 9908 7328 10007
rect 8754 10004 8760 10016
rect 8812 10004 8818 10056
rect 9140 10044 9168 10075
rect 9398 10072 9404 10124
rect 9456 10112 9462 10124
rect 10965 10115 11023 10121
rect 10965 10112 10977 10115
rect 9456 10084 10977 10112
rect 9456 10072 9462 10084
rect 10965 10081 10977 10084
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 11146 10072 11152 10124
rect 11204 10072 11210 10124
rect 11422 10072 11428 10124
rect 11480 10072 11486 10124
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 12268 10121 12296 10152
rect 12710 10140 12716 10152
rect 12768 10140 12774 10192
rect 13740 10180 13768 10220
rect 12912 10152 13400 10180
rect 12912 10121 12940 10152
rect 12253 10115 12311 10121
rect 12253 10112 12265 10115
rect 11572 10084 12265 10112
rect 11572 10072 11578 10084
rect 12253 10081 12265 10084
rect 12299 10081 12311 10115
rect 12253 10075 12311 10081
rect 12345 10115 12403 10121
rect 12345 10081 12357 10115
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10081 12495 10115
rect 12437 10075 12495 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 12667 10084 12909 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 11057 10047 11115 10053
rect 11057 10044 11069 10047
rect 9140 10016 11069 10044
rect 11057 10013 11069 10016
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 12066 10004 12072 10056
rect 12124 10044 12130 10056
rect 12360 10044 12388 10075
rect 12124 10016 12388 10044
rect 12124 10004 12130 10016
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 9033 9979 9091 9985
rect 9033 9976 9045 9979
rect 8076 9948 9045 9976
rect 8076 9936 8082 9948
rect 9033 9945 9045 9948
rect 9079 9945 9091 9979
rect 12452 9976 12480 10075
rect 13078 10072 13084 10124
rect 13136 10072 13142 10124
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 13262 10004 13268 10056
rect 13320 10004 13326 10056
rect 13372 10044 13400 10152
rect 13464 10152 13768 10180
rect 15013 10183 15071 10189
rect 13464 10124 13492 10152
rect 15013 10149 15025 10183
rect 15059 10149 15071 10183
rect 15013 10143 15071 10149
rect 13446 10072 13452 10124
rect 13504 10072 13510 10124
rect 13722 10072 13728 10124
rect 13780 10072 13786 10124
rect 14090 10112 14096 10124
rect 13832 10084 14096 10112
rect 13832 10044 13860 10084
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 14826 10121 14832 10124
rect 14824 10075 14832 10121
rect 14826 10072 14832 10075
rect 14884 10072 14890 10124
rect 14921 10115 14979 10121
rect 14921 10081 14933 10115
rect 14967 10081 14979 10115
rect 14921 10075 14979 10081
rect 13372 10016 13860 10044
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14001 10047 14059 10053
rect 14001 10044 14013 10047
rect 13964 10016 14013 10044
rect 13964 10004 13970 10016
rect 14001 10013 14013 10016
rect 14047 10044 14059 10047
rect 14366 10044 14372 10056
rect 14047 10016 14372 10044
rect 14047 10013 14059 10016
rect 14001 10007 14059 10013
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14936 10044 14964 10075
rect 14844 10016 14964 10044
rect 14645 9979 14703 9985
rect 14645 9976 14657 9979
rect 12452 9948 14657 9976
rect 9033 9939 9091 9945
rect 14645 9945 14657 9948
rect 14691 9945 14703 9979
rect 14645 9939 14703 9945
rect 6880 9880 7328 9908
rect 6880 9868 6886 9880
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13722 9908 13728 9920
rect 13228 9880 13728 9908
rect 13228 9868 13234 9880
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 13814 9868 13820 9920
rect 13872 9868 13878 9920
rect 13909 9911 13967 9917
rect 13909 9877 13921 9911
rect 13955 9908 13967 9911
rect 13998 9908 14004 9920
rect 13955 9880 14004 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 13998 9868 14004 9880
rect 14056 9868 14062 9920
rect 14844 9908 14872 10016
rect 15028 9976 15056 10143
rect 15194 10072 15200 10124
rect 15252 10072 15258 10124
rect 15304 10121 15332 10220
rect 16206 10208 16212 10260
rect 16264 10208 16270 10260
rect 15470 10140 15476 10192
rect 15528 10180 15534 10192
rect 15528 10152 16344 10180
rect 15528 10140 15534 10152
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 15378 10072 15384 10124
rect 15436 10072 15442 10124
rect 15562 10072 15568 10124
rect 15620 10072 15626 10124
rect 16114 10072 16120 10124
rect 16172 10072 16178 10124
rect 16316 10121 16344 10152
rect 16301 10115 16359 10121
rect 16301 10081 16313 10115
rect 16347 10112 16359 10115
rect 16482 10112 16488 10124
rect 16347 10084 16488 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 15028 9948 15393 9976
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 15562 9908 15568 9920
rect 14844 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 4617 9707 4675 9713
rect 4617 9704 4629 9707
rect 4580 9676 4629 9704
rect 4580 9664 4586 9676
rect 4617 9673 4629 9676
rect 4663 9673 4675 9707
rect 4617 9667 4675 9673
rect 5626 9664 5632 9716
rect 5684 9664 5690 9716
rect 6362 9664 6368 9716
rect 6420 9664 6426 9716
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6512 9676 6745 9704
rect 6512 9664 6518 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 11146 9664 11152 9716
rect 11204 9664 11210 9716
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 12124 9676 12173 9704
rect 12124 9664 12130 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 13081 9707 13139 9713
rect 13081 9704 13093 9707
rect 12492 9676 13093 9704
rect 12492 9664 12498 9676
rect 13081 9673 13093 9676
rect 13127 9704 13139 9707
rect 13170 9704 13176 9716
rect 13127 9676 13176 9704
rect 13127 9673 13139 9676
rect 13081 9667 13139 9673
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13262 9664 13268 9716
rect 13320 9704 13326 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 13320 9676 13553 9704
rect 13320 9664 13326 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 15105 9707 15163 9713
rect 15105 9704 15117 9707
rect 14884 9676 15117 9704
rect 14884 9664 14890 9676
rect 15105 9673 15117 9676
rect 15151 9673 15163 9707
rect 15105 9667 15163 9673
rect 5442 9636 5448 9648
rect 4632 9608 5448 9636
rect 4632 9500 4660 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 4706 9528 4712 9580
rect 4764 9568 4770 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4764 9540 4905 9568
rect 4764 9528 4770 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5644 9568 5672 9664
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6319 9608 6653 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7285 9639 7343 9645
rect 7285 9636 7297 9639
rect 6972 9608 7297 9636
rect 6972 9596 6978 9608
rect 7285 9605 7297 9608
rect 7331 9636 7343 9639
rect 8202 9636 8208 9648
rect 7331 9608 8208 9636
rect 7331 9605 7343 9608
rect 7285 9599 7343 9605
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 9769 9639 9827 9645
rect 9769 9636 9781 9639
rect 9732 9608 9781 9636
rect 9732 9596 9738 9608
rect 9769 9605 9781 9608
rect 9815 9605 9827 9639
rect 9769 9599 9827 9605
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 13446 9636 13452 9648
rect 11664 9608 13124 9636
rect 11664 9596 11670 9608
rect 5132 9540 5672 9568
rect 6457 9571 6515 9577
rect 5132 9528 5138 9540
rect 6457 9537 6469 9571
rect 6503 9537 6515 9571
rect 6457 9531 6515 9537
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4632 9472 4813 9500
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 5000 9432 5028 9463
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 5868 9472 6193 9500
rect 5868 9460 5874 9472
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6472 9432 6500 9531
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6788 9540 6960 9568
rect 6788 9528 6794 9540
rect 6822 9460 6828 9512
rect 6880 9460 6886 9512
rect 6932 9500 6960 9540
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 7064 9540 7113 9568
rect 7064 9528 7070 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 8018 9568 8024 9580
rect 7101 9531 7159 9537
rect 7484 9540 8024 9568
rect 7484 9509 7512 9540
rect 8018 9528 8024 9540
rect 8076 9528 8082 9580
rect 9398 9568 9404 9580
rect 8956 9540 9404 9568
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 6932 9472 7389 9500
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 7650 9460 7656 9512
rect 7708 9460 7714 9512
rect 8956 9509 8984 9540
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11563 9540 12112 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 7561 9435 7619 9441
rect 7561 9432 7573 9435
rect 4396 9404 6040 9432
rect 6472 9404 7573 9432
rect 4396 9392 4402 9404
rect 6012 9376 6040 9404
rect 7561 9401 7573 9404
rect 7607 9401 7619 9435
rect 9140 9432 9168 9463
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 11054 9460 11060 9512
rect 11112 9460 11118 9512
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9469 11391 9503
rect 11333 9463 11391 9469
rect 11425 9503 11483 9509
rect 11425 9469 11437 9503
rect 11471 9469 11483 9503
rect 11425 9463 11483 9469
rect 9490 9432 9496 9444
rect 9140 9404 9496 9432
rect 7561 9395 7619 9401
rect 9490 9392 9496 9404
rect 9548 9432 9554 9444
rect 10870 9432 10876 9444
rect 9548 9404 10876 9432
rect 9548 9392 9554 9404
rect 10870 9392 10876 9404
rect 10928 9432 10934 9444
rect 11348 9432 11376 9463
rect 10928 9404 11376 9432
rect 11440 9432 11468 9463
rect 11606 9460 11612 9512
rect 11664 9460 11670 9512
rect 12084 9500 12112 9540
rect 12250 9528 12256 9580
rect 12308 9568 12314 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12308 9540 12541 9568
rect 12308 9528 12314 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12986 9568 12992 9580
rect 12676 9540 12992 9568
rect 12676 9528 12682 9540
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13096 9568 13124 9608
rect 13372 9608 13452 9636
rect 13372 9568 13400 9608
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15654 9636 15660 9648
rect 15252 9608 15660 9636
rect 15252 9596 15258 9608
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 15838 9596 15844 9648
rect 15896 9596 15902 9648
rect 16577 9639 16635 9645
rect 16577 9605 16589 9639
rect 16623 9605 16635 9639
rect 16577 9599 16635 9605
rect 15212 9568 15240 9596
rect 16022 9568 16028 9580
rect 13096 9540 13400 9568
rect 13648 9540 14964 9568
rect 15212 9540 15333 9568
rect 12342 9509 12348 9512
rect 12341 9500 12348 9509
rect 12084 9472 12348 9500
rect 12341 9463 12348 9472
rect 12342 9460 12348 9463
rect 12400 9460 12406 9512
rect 12434 9460 12440 9512
rect 12492 9460 12498 9512
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 13096 9509 13124 9540
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 12066 9432 12072 9444
rect 11440 9404 12072 9432
rect 10928 9392 10934 9404
rect 12066 9392 12072 9404
rect 12124 9392 12130 9444
rect 12912 9432 12940 9463
rect 13648 9432 13676 9540
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 12728 9404 13676 9432
rect 12728 9376 12756 9404
rect 13832 9376 13860 9463
rect 13998 9460 14004 9512
rect 14056 9509 14062 9512
rect 14056 9503 14085 9509
rect 14073 9469 14085 9503
rect 14056 9463 14085 9469
rect 14056 9460 14062 9463
rect 14182 9460 14188 9512
rect 14240 9460 14246 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 14936 9509 14964 9540
rect 14645 9503 14703 9509
rect 14645 9500 14657 9503
rect 14516 9472 14657 9500
rect 14516 9460 14522 9472
rect 14645 9469 14657 9472
rect 14691 9469 14703 9503
rect 14645 9463 14703 9469
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9432 13967 9435
rect 14366 9432 14372 9444
rect 13955 9404 14372 9432
rect 13955 9401 13967 9404
rect 13909 9395 13967 9401
rect 14366 9392 14372 9404
rect 14424 9392 14430 9444
rect 14936 9432 14964 9463
rect 15194 9460 15200 9512
rect 15252 9460 15258 9512
rect 15305 9509 15333 9540
rect 15488 9540 16028 9568
rect 15488 9509 15516 9540
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 16592 9568 16620 9599
rect 16316 9540 16620 9568
rect 15290 9503 15348 9509
rect 15290 9469 15302 9503
rect 15336 9469 15348 9503
rect 15290 9463 15348 9469
rect 15473 9503 15531 9509
rect 15473 9469 15485 9503
rect 15519 9469 15531 9503
rect 15473 9463 15531 9469
rect 15703 9503 15761 9509
rect 15703 9469 15715 9503
rect 15749 9500 15761 9503
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15749 9472 15945 9500
rect 15749 9469 15761 9472
rect 15703 9463 15761 9469
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 16206 9460 16212 9512
rect 16264 9460 16270 9512
rect 14936 9404 15516 9432
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 6270 9364 6276 9376
rect 6052 9336 6276 9364
rect 6052 9324 6058 9336
rect 6270 9324 6276 9336
rect 6328 9364 6334 9376
rect 6546 9364 6552 9376
rect 6328 9336 6552 9364
rect 6328 9324 6334 9336
rect 6546 9324 6552 9336
rect 6604 9364 6610 9376
rect 7006 9364 7012 9376
rect 6604 9336 7012 9364
rect 6604 9324 6610 9336
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 7742 9324 7748 9376
rect 7800 9364 7806 9376
rect 8570 9364 8576 9376
rect 7800 9336 8576 9364
rect 7800 9324 7806 9336
rect 8570 9324 8576 9336
rect 8628 9364 8634 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8628 9336 8769 9364
rect 8628 9324 8634 9336
rect 8757 9333 8769 9336
rect 8803 9364 8815 9367
rect 9030 9364 9036 9376
rect 8803 9336 9036 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10962 9364 10968 9376
rect 10560 9336 10968 9364
rect 10560 9324 10566 9336
rect 10962 9324 10968 9336
rect 11020 9364 11026 9376
rect 12434 9364 12440 9376
rect 11020 9336 12440 9364
rect 11020 9324 11026 9336
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13136 9336 13277 9364
rect 13136 9324 13142 9336
rect 13265 9333 13277 9336
rect 13311 9364 13323 9367
rect 13630 9364 13636 9376
rect 13311 9336 13636 9364
rect 13311 9333 13323 9336
rect 13265 9327 13323 9333
rect 13630 9324 13636 9336
rect 13688 9324 13694 9376
rect 13814 9324 13820 9376
rect 13872 9324 13878 9376
rect 13998 9324 14004 9376
rect 14056 9364 14062 9376
rect 14737 9367 14795 9373
rect 14737 9364 14749 9367
rect 14056 9336 14749 9364
rect 14056 9324 14062 9336
rect 14737 9333 14749 9336
rect 14783 9364 14795 9367
rect 15378 9364 15384 9376
rect 14783 9336 15384 9364
rect 14783 9333 14795 9336
rect 14737 9327 14795 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15488 9364 15516 9404
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 16316 9432 16344 9540
rect 16390 9460 16396 9512
rect 16448 9460 16454 9512
rect 16482 9460 16488 9512
rect 16540 9460 16546 9512
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16684 9472 16865 9500
rect 15620 9404 16344 9432
rect 15620 9392 15626 9404
rect 16574 9392 16580 9444
rect 16632 9392 16638 9444
rect 15930 9364 15936 9376
rect 15488 9336 15936 9364
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16390 9324 16396 9376
rect 16448 9364 16454 9376
rect 16684 9364 16712 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 16448 9336 16712 9364
rect 16448 9324 16454 9336
rect 16758 9324 16764 9376
rect 16816 9324 16822 9376
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 6748 9132 7052 9160
rect 6748 9101 6776 9132
rect 6733 9095 6791 9101
rect 6733 9061 6745 9095
rect 6779 9061 6791 9095
rect 6733 9055 6791 9061
rect 6822 9052 6828 9104
rect 6880 9092 6886 9104
rect 6933 9095 6991 9101
rect 6933 9092 6945 9095
rect 6880 9064 6945 9092
rect 6880 9052 6886 9064
rect 6932 9061 6945 9064
rect 6979 9061 6991 9095
rect 7024 9092 7052 9132
rect 7098 9120 7104 9172
rect 7156 9120 7162 9172
rect 7650 9120 7656 9172
rect 7708 9160 7714 9172
rect 8110 9160 8116 9172
rect 7708 9132 8116 9160
rect 7708 9120 7714 9132
rect 8110 9120 8116 9132
rect 8168 9160 8174 9172
rect 8849 9163 8907 9169
rect 8849 9160 8861 9163
rect 8168 9132 8861 9160
rect 8168 9120 8174 9132
rect 8849 9129 8861 9132
rect 8895 9129 8907 9163
rect 8849 9123 8907 9129
rect 8956 9132 9260 9160
rect 7282 9092 7288 9104
rect 7024 9064 7288 9092
rect 6932 9055 6991 9061
rect 6546 8984 6552 9036
rect 6604 9024 6610 9036
rect 6932 9024 6960 9055
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 7742 9092 7748 9104
rect 7392 9064 7748 9092
rect 7392 9033 7420 9064
rect 7742 9052 7748 9064
rect 7800 9092 7806 9104
rect 8021 9095 8079 9101
rect 8021 9092 8033 9095
rect 7800 9064 8033 9092
rect 7800 9052 7806 9064
rect 8021 9061 8033 9064
rect 8067 9061 8079 9095
rect 8021 9055 8079 9061
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9061 8539 9095
rect 8481 9055 8539 9061
rect 6604 8996 6960 9024
rect 6604 8984 6610 8996
rect 6932 8888 6960 8996
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 7558 8984 7564 9036
rect 7616 8984 7622 9036
rect 7834 8984 7840 9036
rect 7892 8984 7898 9036
rect 8343 9027 8401 9033
rect 8343 9024 8355 9027
rect 8097 9017 8155 9023
rect 8097 9014 8109 9017
rect 8036 8986 8109 9014
rect 7576 8956 7604 8984
rect 8036 8956 8064 8986
rect 8097 8983 8109 8986
rect 8143 8983 8155 9017
rect 8097 8977 8155 8983
rect 8220 8996 8355 9024
rect 7576 8928 8064 8956
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 6932 8860 7665 8888
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 7926 8848 7932 8900
rect 7984 8888 7990 8900
rect 8220 8888 8248 8996
rect 8343 8993 8355 8996
rect 8389 8993 8401 9027
rect 8496 9022 8524 9055
rect 8570 9052 8576 9104
rect 8628 9052 8634 9104
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 8956 9092 8984 9132
rect 8720 9064 8984 9092
rect 9017 9095 9075 9101
rect 8720 9052 8726 9064
rect 9017 9061 9029 9095
rect 9063 9092 9075 9095
rect 9122 9092 9128 9104
rect 9063 9064 9128 9092
rect 9063 9061 9075 9064
rect 9017 9055 9075 9061
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9232 9101 9260 9132
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10318 9160 10324 9172
rect 10192 9132 10324 9160
rect 10192 9120 10198 9132
rect 10318 9120 10324 9132
rect 10376 9120 10382 9172
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11422 9160 11428 9172
rect 11379 9132 11428 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 12710 9160 12716 9172
rect 12452 9132 12716 9160
rect 9217 9095 9275 9101
rect 9217 9061 9229 9095
rect 9263 9061 9275 9095
rect 9861 9095 9919 9101
rect 9861 9092 9873 9095
rect 9217 9055 9275 9061
rect 9324 9064 9873 9092
rect 8588 9022 8708 9024
rect 8496 8996 8708 9022
rect 8496 8994 8616 8996
rect 8343 8987 8401 8993
rect 8680 8968 8708 8996
rect 8754 8984 8760 9036
rect 8812 9024 8818 9036
rect 9324 9024 9352 9064
rect 9861 9061 9873 9064
rect 9907 9061 9919 9095
rect 9861 9055 9919 9061
rect 8812 8996 9352 9024
rect 8812 8984 8818 8996
rect 9490 8984 9496 9036
rect 9548 8984 9554 9036
rect 9582 8984 9588 9036
rect 9640 8984 9646 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 8662 8916 8668 8968
rect 8720 8916 8726 8968
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9214 8956 9220 8968
rect 8996 8928 9220 8956
rect 8996 8916 9002 8928
rect 7984 8860 8248 8888
rect 9140 8888 9168 8928
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9692 8956 9720 8987
rect 9766 8984 9772 9036
rect 9824 8984 9830 9036
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10962 9024 10968 9036
rect 9999 8996 10968 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10962 8984 10968 8996
rect 11020 9024 11026 9036
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 11020 8996 11161 9024
rect 11020 8984 11026 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 11514 8984 11520 9036
rect 11572 8984 11578 9036
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 11974 9024 11980 9036
rect 11839 8996 11980 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 11974 8984 11980 8996
rect 12032 9024 12038 9036
rect 12452 9024 12480 9132
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 13081 9163 13139 9169
rect 13081 9129 13093 9163
rect 13127 9160 13139 9163
rect 13725 9163 13783 9169
rect 13127 9132 13676 9160
rect 13127 9129 13139 9132
rect 13081 9123 13139 9129
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12032 8996 12541 9024
rect 12032 8984 12038 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 12618 8984 12624 9036
rect 12676 8984 12682 9036
rect 12713 9027 12771 9033
rect 12713 8993 12725 9027
rect 12759 8993 12771 9027
rect 12713 8987 12771 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 8993 12955 9027
rect 12897 8987 12955 8993
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 10226 8956 10232 8968
rect 9692 8928 10232 8956
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12728 8956 12756 8987
rect 12492 8928 12756 8956
rect 12912 8956 12940 8987
rect 12986 8956 12992 8968
rect 12912 8928 12992 8956
rect 12492 8916 12498 8928
rect 9140 8860 9812 8888
rect 7984 8848 7990 8860
rect 9784 8832 9812 8860
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10410 8888 10416 8900
rect 10008 8860 10416 8888
rect 10008 8848 10014 8860
rect 10410 8848 10416 8860
rect 10468 8848 10474 8900
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 11112 8860 11652 8888
rect 11112 8848 11118 8860
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 5902 8820 5908 8832
rect 5500 8792 5908 8820
rect 5500 8780 5506 8792
rect 5902 8780 5908 8792
rect 5960 8820 5966 8832
rect 6914 8820 6920 8832
rect 5960 8792 6920 8820
rect 5960 8780 5966 8792
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7432 8792 7481 8820
rect 7432 8780 7438 8792
rect 7469 8789 7481 8792
rect 7515 8820 7527 8823
rect 8018 8820 8024 8832
rect 7515 8792 8024 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8202 8780 8208 8832
rect 8260 8780 8266 8832
rect 9030 8829 9036 8832
rect 9011 8823 9036 8829
rect 9011 8789 9023 8823
rect 9011 8783 9036 8789
rect 9030 8780 9036 8783
rect 9088 8780 9094 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 11238 8820 11244 8832
rect 9824 8792 11244 8820
rect 9824 8780 9830 8792
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11624 8829 11652 8860
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 12618 8820 12624 8832
rect 11655 8792 12624 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 12728 8820 12756 8928
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 13096 8956 13124 8987
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13262 8984 13268 9036
rect 13320 8984 13326 9036
rect 13446 8984 13452 9036
rect 13504 8984 13510 9036
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13648 9024 13676 9132
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 14182 9160 14188 9172
rect 13771 9132 14188 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 14366 9120 14372 9172
rect 14424 9160 14430 9172
rect 16574 9160 16580 9172
rect 14424 9132 16580 9160
rect 14424 9120 14430 9132
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 13722 9024 13728 9036
rect 13648 8996 13728 9024
rect 13541 8987 13599 8993
rect 13354 8956 13360 8968
rect 13096 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8956 13418 8968
rect 13556 8956 13584 8987
rect 13722 8984 13728 8996
rect 13780 9024 13786 9036
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13780 8996 13829 9024
rect 13780 8984 13786 8996
rect 13817 8993 13829 8996
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 14090 8984 14096 9036
rect 14148 9024 14154 9036
rect 14918 9024 14924 9036
rect 14148 8996 14924 9024
rect 14148 8984 14154 8996
rect 14918 8984 14924 8996
rect 14976 8984 14982 9036
rect 15378 8984 15384 9036
rect 15436 8984 15442 9036
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 8993 15623 9027
rect 15565 8987 15623 8993
rect 13412 8928 13584 8956
rect 13412 8916 13418 8928
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 13688 8928 13921 8956
rect 13688 8916 13694 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 13909 8919 13967 8925
rect 15010 8916 15016 8968
rect 15068 8956 15074 8968
rect 15580 8956 15608 8987
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16264 8996 16497 9024
rect 16264 8984 16270 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 15068 8928 15608 8956
rect 15068 8916 15074 8928
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15988 8928 16313 8956
rect 15988 8916 15994 8928
rect 16301 8925 16313 8928
rect 16347 8925 16359 8959
rect 16500 8956 16528 8987
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16632 8996 16957 9024
rect 16632 8984 16638 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 16945 8987 17003 8993
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 9024 17187 9027
rect 17218 9024 17224 9036
rect 17175 8996 17224 9024
rect 17175 8993 17187 8996
rect 17129 8987 17187 8993
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 16500 8928 16620 8956
rect 16301 8919 16359 8925
rect 13004 8888 13032 8916
rect 16592 8900 16620 8928
rect 14458 8888 14464 8900
rect 13004 8860 14464 8888
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 16574 8848 16580 8900
rect 16632 8848 16638 8900
rect 13078 8820 13084 8832
rect 12728 8792 13084 8820
rect 13078 8780 13084 8792
rect 13136 8820 13142 8832
rect 13814 8820 13820 8832
rect 13136 8792 13820 8820
rect 13136 8780 13142 8792
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14274 8780 14280 8832
rect 14332 8780 14338 8832
rect 15381 8823 15439 8829
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 15562 8820 15568 8832
rect 15427 8792 15568 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16390 8820 16396 8832
rect 16172 8792 16396 8820
rect 16172 8780 16178 8792
rect 16390 8780 16396 8792
rect 16448 8820 16454 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16448 8792 16681 8820
rect 16448 8780 16454 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 16758 8780 16764 8832
rect 16816 8780 16822 8832
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 4614 8616 4620 8628
rect 4295 8588 4620 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 9180 8588 9413 8616
rect 9180 8576 9186 8588
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 10134 8576 10140 8628
rect 10192 8616 10198 8628
rect 10594 8616 10600 8628
rect 10192 8588 10600 8616
rect 10192 8576 10198 8588
rect 10594 8576 10600 8588
rect 10652 8616 10658 8628
rect 11422 8616 11428 8628
rect 10652 8588 11428 8616
rect 10652 8576 10658 8588
rect 11422 8576 11428 8588
rect 11480 8576 11486 8628
rect 13538 8576 13544 8628
rect 13596 8576 13602 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 13648 8588 14841 8616
rect 3605 8551 3663 8557
rect 3605 8517 3617 8551
rect 3651 8548 3663 8551
rect 4062 8548 4068 8560
rect 3651 8520 4068 8548
rect 3651 8517 3663 8520
rect 3605 8511 3663 8517
rect 4062 8508 4068 8520
rect 4120 8548 4126 8560
rect 9217 8551 9275 8557
rect 4120 8520 4476 8548
rect 4120 8508 4126 8520
rect 4448 8489 4476 8520
rect 5184 8520 6408 8548
rect 4433 8483 4491 8489
rect 3988 8452 4384 8480
rect 3786 8372 3792 8424
rect 3844 8372 3850 8424
rect 3988 8421 4016 8452
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4246 8372 4252 8424
rect 4304 8372 4310 8424
rect 4356 8412 4384 8452
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4801 8483 4859 8489
rect 4801 8480 4813 8483
rect 4580 8452 4813 8480
rect 4580 8440 4586 8452
rect 4632 8421 4660 8452
rect 4801 8449 4813 8452
rect 4847 8449 4859 8483
rect 4982 8480 4988 8492
rect 4801 8443 4859 8449
rect 4908 8452 4988 8480
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4356 8384 4629 8412
rect 4617 8381 4629 8384
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 4908 8421 4936 8452
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5184 8421 5212 8520
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 6380 8480 6408 8520
rect 9217 8517 9229 8551
rect 9263 8517 9275 8551
rect 9508 8548 9536 8576
rect 9766 8548 9772 8560
rect 9217 8511 9275 8517
rect 9416 8520 9536 8548
rect 9646 8520 9772 8548
rect 6730 8480 6736 8492
rect 5491 8452 6132 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 6104 8424 6132 8452
rect 6380 8452 6736 8480
rect 4893 8415 4951 8421
rect 4893 8381 4905 8415
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5997 8415 6055 8421
rect 5997 8412 6009 8415
rect 5583 8384 6009 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5997 8381 6009 8384
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4525 8347 4583 8353
rect 4525 8344 4537 8347
rect 3927 8316 4537 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4525 8313 4537 8316
rect 4571 8344 4583 8347
rect 4985 8347 5043 8353
rect 4985 8344 4997 8347
rect 4571 8316 4997 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 4985 8313 4997 8316
rect 5031 8313 5043 8347
rect 4985 8307 5043 8313
rect 5276 8344 5304 8375
rect 5626 8344 5632 8356
rect 5276 8316 5632 8344
rect 4154 8236 4160 8288
rect 4212 8236 4218 8288
rect 4706 8236 4712 8288
rect 4764 8276 4770 8288
rect 5276 8276 5304 8316
rect 5626 8304 5632 8316
rect 5684 8304 5690 8356
rect 6012 8344 6040 8375
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6181 8415 6239 8421
rect 6181 8412 6193 8415
rect 6144 8384 6193 8412
rect 6144 8372 6150 8384
rect 6181 8381 6193 8384
rect 6227 8381 6239 8415
rect 6181 8375 6239 8381
rect 6270 8372 6276 8424
rect 6328 8372 6334 8424
rect 6380 8421 6408 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7834 8480 7840 8492
rect 7024 8452 7840 8480
rect 7024 8424 7052 8452
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 9232 8480 9260 8511
rect 8772 8452 9260 8480
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6454 8412 6460 8424
rect 6411 8384 6460 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 6546 8372 6552 8424
rect 6604 8372 6610 8424
rect 6917 8415 6975 8421
rect 6917 8381 6929 8415
rect 6963 8412 6975 8415
rect 7006 8412 7012 8424
rect 6963 8384 7012 8412
rect 6963 8381 6975 8384
rect 6917 8375 6975 8381
rect 7006 8372 7012 8384
rect 7064 8372 7070 8424
rect 7190 8372 7196 8424
rect 7248 8412 7254 8424
rect 7926 8412 7932 8424
rect 7248 8384 7932 8412
rect 7248 8372 7254 8384
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8772 8421 8800 8452
rect 8757 8415 8815 8421
rect 8757 8381 8769 8415
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8849 8415 8907 8421
rect 8849 8381 8861 8415
rect 8895 8412 8907 8415
rect 9416 8412 9444 8520
rect 9493 8483 9551 8489
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 9646 8480 9674 8520
rect 9766 8508 9772 8520
rect 9824 8548 9830 8560
rect 9950 8548 9956 8560
rect 9824 8520 9956 8548
rect 9824 8508 9830 8520
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10502 8548 10508 8560
rect 10428 8520 10508 8548
rect 9539 8452 9674 8480
rect 9861 8483 9919 8489
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 9861 8449 9873 8483
rect 9907 8480 9919 8483
rect 10134 8480 10140 8492
rect 9907 8452 10140 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8480 10379 8483
rect 10428 8480 10456 8520
rect 10502 8508 10508 8520
rect 10560 8508 10566 8560
rect 10870 8508 10876 8560
rect 10928 8508 10934 8560
rect 10962 8508 10968 8560
rect 11020 8508 11026 8560
rect 12618 8508 12624 8560
rect 12676 8548 12682 8560
rect 13446 8548 13452 8560
rect 12676 8520 13452 8548
rect 12676 8508 12682 8520
rect 13446 8508 13452 8520
rect 13504 8548 13510 8560
rect 13648 8548 13676 8588
rect 14829 8585 14841 8588
rect 14875 8616 14887 8619
rect 14918 8616 14924 8628
rect 14875 8588 14924 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 14918 8576 14924 8588
rect 14976 8576 14982 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 16206 8616 16212 8628
rect 15620 8588 16212 8616
rect 15620 8576 15626 8588
rect 16206 8576 16212 8588
rect 16264 8616 16270 8628
rect 17218 8616 17224 8628
rect 16264 8588 17224 8616
rect 16264 8576 16270 8588
rect 17218 8576 17224 8588
rect 17276 8576 17282 8628
rect 14274 8548 14280 8560
rect 13504 8520 13676 8548
rect 13740 8520 14280 8548
rect 13504 8508 13510 8520
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 10367 8452 10456 8480
rect 11716 8452 11989 8480
rect 10367 8449 10379 8452
rect 10321 8443 10379 8449
rect 8895 8384 9444 8412
rect 8895 8381 8907 8384
rect 8849 8375 8907 8381
rect 9582 8372 9588 8424
rect 9640 8372 9646 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9950 8412 9956 8424
rect 9723 8384 9956 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10045 8415 10103 8421
rect 10045 8381 10057 8415
rect 10091 8412 10103 8415
rect 10410 8412 10416 8424
rect 10091 8384 10416 8412
rect 10091 8381 10103 8384
rect 10045 8375 10103 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10594 8378 10600 8424
rect 10520 8372 10600 8378
rect 10652 8372 10658 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 10735 8384 11621 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6012 8316 6837 8344
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 8938 8304 8944 8356
rect 8996 8304 9002 8356
rect 9125 8347 9183 8353
rect 9125 8313 9137 8347
rect 9171 8344 9183 8347
rect 9490 8344 9496 8356
rect 9171 8316 9496 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10226 8344 10232 8356
rect 9784 8316 10232 8344
rect 4764 8248 5304 8276
rect 5644 8276 5672 8304
rect 6270 8276 6276 8288
rect 5644 8248 6276 8276
rect 4764 8236 4770 8248
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 7098 8236 7104 8288
rect 7156 8236 7162 8288
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 9784 8285 9812 8316
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10520 8350 10640 8372
rect 8573 8279 8631 8285
rect 8573 8276 8585 8279
rect 8352 8248 8585 8276
rect 8352 8236 8358 8248
rect 8573 8245 8585 8248
rect 8619 8245 8631 8279
rect 8573 8239 8631 8245
rect 9769 8279 9827 8285
rect 9769 8245 9781 8279
rect 9815 8245 9827 8279
rect 9769 8239 9827 8245
rect 9953 8279 10011 8285
rect 9953 8245 9965 8279
rect 9999 8276 10011 8279
rect 10042 8276 10048 8288
rect 9999 8248 10048 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 10520 8285 10548 8350
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 11149 8347 11207 8353
rect 11149 8344 11161 8347
rect 11112 8316 11161 8344
rect 11112 8304 11118 8316
rect 11149 8313 11161 8316
rect 11195 8313 11207 8347
rect 11149 8307 11207 8313
rect 11333 8347 11391 8353
rect 11333 8313 11345 8347
rect 11379 8344 11391 8347
rect 11422 8344 11428 8356
rect 11379 8316 11428 8344
rect 11379 8313 11391 8316
rect 11333 8307 11391 8313
rect 11422 8304 11428 8316
rect 11480 8304 11486 8356
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8344 11575 8347
rect 11716 8344 11744 8452
rect 11977 8449 11989 8452
rect 12023 8480 12035 8483
rect 13262 8480 13268 8492
rect 12023 8452 13268 8480
rect 12023 8449 12035 8452
rect 11977 8443 12035 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 11882 8412 11888 8424
rect 11839 8384 11888 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 13740 8421 13768 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 14461 8551 14519 8557
rect 14461 8517 14473 8551
rect 14507 8517 14519 8551
rect 14461 8511 14519 8517
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8517 15991 8551
rect 15933 8511 15991 8517
rect 14476 8480 14504 8511
rect 15948 8480 15976 8511
rect 13832 8452 14504 8480
rect 14844 8452 15976 8480
rect 13832 8421 13860 8452
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8381 13875 8415
rect 13817 8375 13875 8381
rect 14182 8372 14188 8424
rect 14240 8372 14246 8424
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14844 8421 14872 8452
rect 16022 8440 16028 8492
rect 16080 8480 16086 8492
rect 16485 8483 16543 8489
rect 16485 8480 16497 8483
rect 16080 8452 16497 8480
rect 16080 8440 16086 8452
rect 16485 8449 16497 8452
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 14645 8415 14703 8421
rect 14645 8412 14657 8415
rect 14332 8384 14657 8412
rect 14332 8372 14338 8384
rect 14645 8381 14657 8384
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 14829 8415 14887 8421
rect 14829 8381 14841 8415
rect 14875 8381 14887 8415
rect 14829 8375 14887 8381
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 15013 8375 15071 8381
rect 15197 8415 15255 8421
rect 15197 8381 15209 8415
rect 15243 8412 15255 8415
rect 15378 8412 15384 8424
rect 15243 8384 15384 8412
rect 15243 8381 15255 8384
rect 15197 8375 15255 8381
rect 11563 8316 11744 8344
rect 11900 8344 11928 8372
rect 11900 8316 13860 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8245 10563 8279
rect 10505 8239 10563 8245
rect 10597 8279 10655 8285
rect 10597 8245 10609 8279
rect 10643 8276 10655 8279
rect 10778 8276 10784 8288
rect 10643 8248 10784 8276
rect 10643 8245 10655 8248
rect 10597 8239 10655 8245
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 10836 8248 11253 8276
rect 10836 8236 10842 8248
rect 11241 8245 11253 8248
rect 11287 8245 11299 8279
rect 11532 8276 11560 8307
rect 11606 8276 11612 8288
rect 11532 8248 11612 8276
rect 11241 8239 11299 8245
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 13832 8276 13860 8316
rect 13906 8304 13912 8356
rect 13964 8304 13970 8356
rect 13998 8304 14004 8356
rect 14056 8353 14062 8356
rect 14056 8347 14085 8353
rect 14073 8313 14085 8347
rect 14458 8344 14464 8356
rect 14056 8307 14085 8313
rect 14200 8316 14464 8344
rect 14056 8304 14062 8307
rect 14200 8276 14228 8316
rect 14458 8304 14464 8316
rect 14516 8344 14522 8356
rect 15028 8344 15056 8375
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 16758 8412 16764 8424
rect 16347 8384 16764 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 16758 8372 16764 8384
rect 16816 8372 16822 8424
rect 14516 8316 15056 8344
rect 14516 8304 14522 8316
rect 16390 8304 16396 8356
rect 16448 8304 16454 8356
rect 13832 8248 14228 8276
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15470 8276 15476 8288
rect 15427 8248 15476 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4246 8072 4252 8084
rect 3927 8044 4252 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 6181 8075 6239 8081
rect 5040 8044 5488 8072
rect 5040 8032 5046 8044
rect 5460 8013 5488 8044
rect 6181 8041 6193 8075
rect 6227 8072 6239 8075
rect 6362 8072 6368 8084
rect 6227 8044 6368 8072
rect 6227 8041 6239 8044
rect 6181 8035 6239 8041
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 6733 8075 6791 8081
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 7190 8072 7196 8084
rect 6779 8044 7196 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 4617 8007 4675 8013
rect 4617 7973 4629 8007
rect 4663 8004 4675 8007
rect 5077 8007 5135 8013
rect 5077 8004 5089 8007
rect 4663 7976 5089 8004
rect 4663 7973 4675 7976
rect 4617 7967 4675 7973
rect 5077 7973 5089 7976
rect 5123 7973 5135 8007
rect 5077 7967 5135 7973
rect 5445 8007 5503 8013
rect 5445 7973 5457 8007
rect 5491 8004 5503 8007
rect 6748 8004 6776 8035
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 10134 8081 10140 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 9640 8044 9965 8072
rect 9640 8032 9646 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 9953 8035 10011 8041
rect 10121 8075 10140 8081
rect 10121 8041 10133 8075
rect 10192 8072 10198 8084
rect 10962 8072 10968 8084
rect 10192 8044 10968 8072
rect 10121 8035 10140 8041
rect 10134 8032 10140 8035
rect 10192 8032 10198 8044
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12032 8044 12909 8072
rect 12032 8032 12038 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 12897 8035 12955 8041
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 13964 8044 15025 8072
rect 13964 8032 13970 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 16206 8032 16212 8084
rect 16264 8072 16270 8084
rect 16758 8072 16764 8084
rect 16264 8044 16764 8072
rect 16264 8032 16270 8044
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 5491 7976 6500 8004
rect 5491 7973 5503 7976
rect 5445 7967 5503 7973
rect 3418 7896 3424 7948
rect 3476 7945 3482 7948
rect 3476 7899 3488 7945
rect 3697 7939 3755 7945
rect 3697 7905 3709 7939
rect 3743 7936 3755 7939
rect 3970 7936 3976 7948
rect 3743 7908 3976 7936
rect 3743 7905 3755 7908
rect 3697 7899 3755 7905
rect 3476 7896 3482 7899
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3844 7840 3893 7868
rect 3844 7828 3850 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 4172 7868 4200 7899
rect 4522 7896 4528 7948
rect 4580 7896 4586 7948
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 4893 7939 4951 7945
rect 4893 7905 4905 7939
rect 4939 7905 4951 7939
rect 4893 7899 4951 7905
rect 4798 7868 4804 7880
rect 4172 7840 4804 7868
rect 3881 7831 3939 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 4908 7868 4936 7899
rect 4982 7896 4988 7948
rect 5040 7896 5046 7948
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5626 7936 5632 7948
rect 5307 7908 5632 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6086 7936 6092 7948
rect 5776 7908 6092 7936
rect 5776 7896 5782 7908
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 6472 7945 6500 7976
rect 6564 7976 6776 8004
rect 6564 7945 6592 7976
rect 9490 7964 9496 8016
rect 9548 8004 9554 8016
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 9548 7976 10333 8004
rect 9548 7964 9554 7976
rect 10321 7973 10333 7976
rect 10367 8004 10379 8007
rect 10870 8004 10876 8016
rect 10367 7976 10876 8004
rect 10367 7973 10379 7976
rect 10321 7967 10379 7973
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 12529 8007 12587 8013
rect 12529 7973 12541 8007
rect 12575 8004 12587 8007
rect 12802 8004 12808 8016
rect 12575 7976 12808 8004
rect 12575 7973 12587 7976
rect 12529 7967 12587 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 13372 8004 13400 8032
rect 16574 8004 16580 8016
rect 13188 7976 13400 8004
rect 15764 7976 16580 8004
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6730 7936 6736 7948
rect 6687 7908 6736 7936
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 6914 7896 6920 7948
rect 6972 7896 6978 7948
rect 9766 7896 9772 7948
rect 9824 7896 9830 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 10134 7936 10140 7948
rect 9907 7908 10140 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 10134 7896 10140 7908
rect 10192 7896 10198 7948
rect 13188 7945 13216 7976
rect 15764 7948 15792 7976
rect 16574 7964 16580 7976
rect 16632 8004 16638 8016
rect 17037 8007 17095 8013
rect 17037 8004 17049 8007
rect 16632 7976 17049 8004
rect 16632 7964 16638 7976
rect 17037 7973 17049 7976
rect 17083 7973 17095 8007
rect 17037 7967 17095 7973
rect 17218 7964 17224 8016
rect 17276 7964 17282 8016
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7905 13231 7939
rect 13173 7899 13231 7905
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7905 13323 7939
rect 13265 7899 13323 7905
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13814 7936 13820 7948
rect 13495 7908 13820 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 4908 7840 5825 7868
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 6656 7840 12434 7868
rect 6656 7800 6684 7840
rect 10226 7800 10232 7812
rect 3988 7772 6684 7800
rect 9876 7772 10232 7800
rect 2317 7735 2375 7741
rect 2317 7701 2329 7735
rect 2363 7732 2375 7735
rect 3988 7732 4016 7772
rect 2363 7704 4016 7732
rect 2363 7701 2375 7704
rect 2317 7695 2375 7701
rect 4062 7692 4068 7744
rect 4120 7692 4126 7744
rect 4338 7692 4344 7744
rect 4396 7692 4402 7744
rect 6638 7692 6644 7744
rect 6696 7732 6702 7744
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 6696 7704 6929 7732
rect 6696 7692 6702 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 6917 7695 6975 7701
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 9876 7741 9904 7772
rect 10226 7760 10232 7772
rect 10284 7760 10290 7812
rect 9493 7735 9551 7741
rect 9493 7732 9505 7735
rect 7984 7704 9505 7732
rect 7984 7692 7990 7704
rect 9493 7701 9505 7704
rect 9539 7701 9551 7735
rect 9493 7695 9551 7701
rect 9861 7735 9919 7741
rect 9861 7701 9873 7735
rect 9907 7701 9919 7735
rect 9861 7695 9919 7701
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10502 7732 10508 7744
rect 10183 7704 10508 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 12406 7732 12434 7840
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 12820 7800 12848 7831
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 13280 7868 13308 7899
rect 13814 7896 13820 7908
rect 13872 7936 13878 7948
rect 15010 7936 15016 7948
rect 13872 7908 15016 7936
rect 13872 7896 13878 7908
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15194 7896 15200 7948
rect 15252 7896 15258 7948
rect 15378 7896 15384 7948
rect 15436 7896 15442 7948
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7905 15531 7939
rect 15473 7899 15531 7905
rect 13538 7868 13544 7880
rect 13280 7840 13544 7868
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 15488 7868 15516 7899
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15620 7908 15669 7936
rect 15620 7896 15626 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 15746 7896 15752 7948
rect 15804 7896 15810 7948
rect 15930 7896 15936 7948
rect 15988 7896 15994 7948
rect 16298 7945 16304 7948
rect 16296 7899 16304 7945
rect 16298 7896 16304 7899
rect 16356 7896 16362 7948
rect 16393 7939 16451 7945
rect 16393 7905 16405 7939
rect 16439 7905 16451 7939
rect 16393 7899 16451 7905
rect 16408 7868 16436 7899
rect 16482 7896 16488 7948
rect 16540 7896 16546 7948
rect 16668 7939 16726 7945
rect 16668 7905 16680 7939
rect 16714 7905 16726 7939
rect 16668 7899 16726 7905
rect 16574 7868 16580 7880
rect 15488 7840 16160 7868
rect 12676 7772 12848 7800
rect 12676 7760 12682 7772
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 16132 7809 16160 7840
rect 16408 7840 16580 7868
rect 16117 7803 16175 7809
rect 14424 7772 16068 7800
rect 14424 7760 14430 7772
rect 13998 7732 14004 7744
rect 12406 7704 14004 7732
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 15930 7692 15936 7744
rect 15988 7692 15994 7744
rect 16040 7732 16068 7772
rect 16117 7769 16129 7803
rect 16163 7769 16175 7803
rect 16117 7763 16175 7769
rect 16408 7732 16436 7840
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 16684 7868 16712 7899
rect 16758 7896 16764 7948
rect 16816 7896 16822 7948
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16684 7840 16865 7868
rect 16776 7812 16804 7840
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 16758 7760 16764 7812
rect 16816 7760 16822 7812
rect 16040 7704 16436 7732
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 3418 7488 3424 7540
rect 3476 7488 3482 7540
rect 3881 7531 3939 7537
rect 3881 7497 3893 7531
rect 3927 7528 3939 7531
rect 4338 7528 4344 7540
rect 3927 7500 4344 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 5074 7488 5080 7540
rect 5132 7488 5138 7540
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6236 7500 6377 7528
rect 6236 7488 6242 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 6512 7500 8064 7528
rect 6512 7488 6518 7500
rect 5442 7460 5448 7472
rect 4908 7432 5448 7460
rect 3602 7284 3608 7336
rect 3660 7284 3666 7336
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7324 3755 7327
rect 3878 7324 3884 7336
rect 3743 7296 3884 7324
rect 3743 7293 3755 7296
rect 3697 7287 3755 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4154 7324 4160 7336
rect 4019 7296 4160 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4798 7284 4804 7336
rect 4856 7284 4862 7336
rect 4908 7333 4936 7432
rect 5442 7420 5448 7432
rect 5500 7460 5506 7472
rect 5902 7460 5908 7472
rect 5500 7432 5908 7460
rect 5500 7420 5506 7432
rect 5902 7420 5908 7432
rect 5960 7420 5966 7472
rect 6730 7420 6736 7472
rect 6788 7460 6794 7472
rect 7466 7460 7472 7472
rect 6788 7432 7472 7460
rect 6788 7420 6794 7432
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 7834 7420 7840 7472
rect 7892 7420 7898 7472
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 7926 7392 7932 7404
rect 5592 7364 5764 7392
rect 5592 7352 5598 7364
rect 5736 7336 5764 7364
rect 7484 7364 7932 7392
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5644 7256 5672 7287
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 5813 7327 5871 7333
rect 5813 7324 5825 7327
rect 5776 7296 5825 7324
rect 5776 7284 5782 7296
rect 5813 7293 5825 7296
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 5960 7296 6377 7324
rect 5960 7284 5966 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7324 6607 7327
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6595 7296 6929 7324
rect 6595 7293 6607 7296
rect 6549 7287 6607 7293
rect 6917 7293 6929 7296
rect 6963 7324 6975 7327
rect 7098 7324 7104 7336
rect 6963 7296 7104 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 6380 7256 6408 7287
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7484 7333 7512 7364
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 7469 7327 7527 7333
rect 7469 7293 7481 7327
rect 7515 7293 7527 7327
rect 7653 7327 7711 7333
rect 7653 7324 7665 7327
rect 7469 7287 7527 7293
rect 7576 7296 7665 7324
rect 7190 7256 7196 7268
rect 5592 7228 5764 7256
rect 6380 7228 7196 7256
rect 5592 7216 5598 7228
rect 5736 7188 5764 7228
rect 7190 7216 7196 7228
rect 7248 7216 7254 7268
rect 6454 7188 6460 7200
rect 5736 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 7098 7148 7104 7200
rect 7156 7188 7162 7200
rect 7576 7188 7604 7296
rect 7653 7293 7665 7296
rect 7699 7293 7711 7327
rect 7653 7287 7711 7293
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7324 7895 7327
rect 8036 7324 8064 7500
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 11333 7531 11391 7537
rect 11333 7497 11345 7531
rect 11379 7528 11391 7531
rect 11974 7528 11980 7540
rect 11379 7500 11980 7528
rect 11379 7497 11391 7500
rect 11333 7491 11391 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12894 7528 12900 7540
rect 12667 7500 12900 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 13688 7500 15301 7528
rect 13688 7488 13694 7500
rect 15289 7497 15301 7500
rect 15335 7528 15347 7531
rect 15746 7528 15752 7540
rect 15335 7500 15752 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 16482 7528 16488 7540
rect 16347 7500 16488 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 16482 7488 16488 7500
rect 16540 7488 16546 7540
rect 12802 7420 12808 7472
rect 12860 7460 12866 7472
rect 13541 7463 13599 7469
rect 13541 7460 13553 7463
rect 12860 7432 13553 7460
rect 12860 7420 12866 7432
rect 13541 7429 13553 7432
rect 13587 7429 13599 7463
rect 13541 7423 13599 7429
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8352 7364 8616 7392
rect 8352 7352 8358 7364
rect 7883 7296 8064 7324
rect 7883 7293 7895 7296
rect 7837 7287 7895 7293
rect 7852 7256 7880 7287
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8588 7333 8616 7364
rect 11514 7352 11520 7404
rect 11572 7392 11578 7404
rect 12345 7395 12403 7401
rect 12345 7392 12357 7395
rect 11572 7364 12357 7392
rect 11572 7352 11578 7364
rect 12345 7361 12357 7364
rect 12391 7361 12403 7395
rect 12345 7355 12403 7361
rect 12986 7352 12992 7404
rect 13044 7392 13050 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 13044 7364 14841 7392
rect 13044 7352 13050 7364
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8260 7296 8401 7324
rect 8260 7284 8266 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 10560 7296 11253 7324
rect 10560 7284 10566 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 12158 7284 12164 7336
rect 12216 7284 12222 7336
rect 12250 7284 12256 7336
rect 12308 7284 12314 7336
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12483 7296 12725 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 13096 7326 13124 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15930 7352 15936 7404
rect 15988 7392 15994 7404
rect 15988 7364 16620 7392
rect 15988 7352 15994 7364
rect 13173 7327 13231 7333
rect 13173 7326 13185 7327
rect 13096 7298 13185 7326
rect 13173 7293 13185 7298
rect 13219 7293 13231 7327
rect 13173 7287 13231 7293
rect 13262 7284 13268 7336
rect 13320 7324 13326 7336
rect 13320 7296 13676 7324
rect 13320 7284 13326 7296
rect 8478 7256 8484 7268
rect 7852 7228 8484 7256
rect 8478 7216 8484 7228
rect 8536 7256 8542 7268
rect 9306 7256 9312 7268
rect 8536 7228 9312 7256
rect 8536 7216 8542 7228
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 12066 7216 12072 7268
rect 12124 7256 12130 7268
rect 13081 7259 13139 7265
rect 13081 7256 13093 7259
rect 12124 7228 13093 7256
rect 12124 7216 12130 7228
rect 13081 7225 13093 7228
rect 13127 7225 13139 7259
rect 13081 7219 13139 7225
rect 13446 7216 13452 7268
rect 13504 7256 13510 7268
rect 13541 7259 13599 7265
rect 13541 7256 13553 7259
rect 13504 7228 13553 7256
rect 13504 7216 13510 7228
rect 13541 7225 13553 7228
rect 13587 7225 13599 7259
rect 13648 7256 13676 7296
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 13872 7296 14473 7324
rect 13872 7284 13878 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 15470 7284 15476 7336
rect 15528 7324 15534 7336
rect 16301 7327 16359 7333
rect 16301 7324 16313 7327
rect 15528 7296 16313 7324
rect 15528 7284 15534 7296
rect 16301 7293 16313 7296
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 16482 7284 16488 7336
rect 16540 7284 16546 7336
rect 16592 7333 16620 7364
rect 16577 7327 16635 7333
rect 16577 7293 16589 7327
rect 16623 7293 16635 7327
rect 16577 7287 16635 7293
rect 16758 7284 16764 7336
rect 16816 7284 16822 7336
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 13648 7228 14657 7256
rect 13541 7219 13599 7225
rect 14645 7225 14657 7228
rect 14691 7256 14703 7259
rect 15194 7256 15200 7268
rect 14691 7228 15200 7256
rect 14691 7225 14703 7228
rect 14645 7219 14703 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 16669 7259 16727 7265
rect 16669 7256 16681 7259
rect 15436 7228 16681 7256
rect 15436 7216 15442 7228
rect 16669 7225 16681 7228
rect 16715 7225 16727 7259
rect 16669 7219 16727 7225
rect 7650 7188 7656 7200
rect 7156 7160 7656 7188
rect 7156 7148 7162 7160
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 12032 7160 13737 7188
rect 12032 7148 12038 7160
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 13725 7151 13783 7157
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 4798 6944 4804 6996
rect 4856 6984 4862 6996
rect 5350 6984 5356 6996
rect 4856 6956 5356 6984
rect 4856 6944 4862 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 6270 6984 6276 6996
rect 5583 6956 6276 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 5552 6916 5580 6947
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 6362 6944 6368 6996
rect 6420 6984 6426 6996
rect 10962 6984 10968 6996
rect 6420 6956 10968 6984
rect 6420 6944 6426 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 12069 6987 12127 6993
rect 12069 6953 12081 6987
rect 12115 6984 12127 6987
rect 12158 6984 12164 6996
rect 12115 6956 12164 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12710 6944 12716 6996
rect 12768 6944 12774 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 15470 6984 15476 6996
rect 12952 6956 15476 6984
rect 12952 6944 12958 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 8202 6916 8208 6928
rect 5276 6888 5580 6916
rect 8036 6888 8208 6916
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 4985 6851 5043 6857
rect 4985 6848 4997 6851
rect 4856 6820 4997 6848
rect 4856 6808 4862 6820
rect 4985 6817 4997 6820
rect 5031 6848 5043 6851
rect 5276 6848 5304 6888
rect 5031 6820 5304 6848
rect 5031 6817 5043 6820
rect 4985 6811 5043 6817
rect 5350 6808 5356 6860
rect 5408 6808 5414 6860
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5491 6820 6040 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5626 6780 5632 6792
rect 5123 6752 5632 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5626 6740 5632 6752
rect 5684 6780 5690 6792
rect 5902 6780 5908 6792
rect 5684 6752 5908 6780
rect 5684 6740 5690 6752
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 4706 6672 4712 6724
rect 4764 6712 4770 6724
rect 6012 6712 6040 6820
rect 7006 6808 7012 6860
rect 7064 6808 7070 6860
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 7466 6808 7472 6860
rect 7524 6808 7530 6860
rect 7650 6808 7656 6860
rect 7708 6808 7714 6860
rect 8036 6857 8064 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 10928 6888 12434 6916
rect 10928 6876 10934 6888
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6817 8079 6851
rect 8021 6811 8079 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8297 6851 8355 6857
rect 8297 6848 8309 6851
rect 8113 6811 8171 6817
rect 8220 6820 8309 6848
rect 7282 6740 7288 6792
rect 7340 6780 7346 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7340 6752 7573 6780
rect 7340 6740 7346 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 8128 6780 8156 6811
rect 8220 6792 8248 6820
rect 8297 6817 8309 6820
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 8829 6851 8887 6857
rect 8829 6848 8841 6851
rect 8720 6820 8841 6848
rect 8720 6808 8726 6820
rect 8829 6817 8841 6820
rect 8875 6817 8887 6851
rect 8829 6811 8887 6817
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 11149 6851 11207 6857
rect 11149 6817 11161 6851
rect 11195 6817 11207 6851
rect 11149 6811 11207 6817
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11471 6820 11560 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 7561 6743 7619 6749
rect 8036 6752 8156 6780
rect 8036 6724 8064 6752
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 7926 6712 7932 6724
rect 4764 6684 7932 6712
rect 4764 6672 4770 6684
rect 7926 6672 7932 6684
rect 7984 6672 7990 6724
rect 8018 6672 8024 6724
rect 8076 6672 8082 6724
rect 9953 6715 10011 6721
rect 9953 6681 9965 6715
rect 9999 6712 10011 6715
rect 10410 6712 10416 6724
rect 9999 6684 10416 6712
rect 9999 6681 10011 6684
rect 9953 6675 10011 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 11164 6712 11192 6811
rect 11422 6712 11428 6724
rect 11164 6684 11428 6712
rect 11422 6672 11428 6684
rect 11480 6672 11486 6724
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4801 6647 4859 6653
rect 4801 6644 4813 6647
rect 4120 6616 4813 6644
rect 4120 6604 4126 6616
rect 4801 6613 4813 6616
rect 4847 6613 4859 6647
rect 4801 6607 4859 6613
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 5169 6647 5227 6653
rect 5169 6644 5181 6647
rect 5132 6616 5181 6644
rect 5132 6604 5138 6616
rect 5169 6613 5181 6616
rect 5215 6613 5227 6647
rect 5169 6607 5227 6613
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5534 6644 5540 6656
rect 5307 6616 5540 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5534 6604 5540 6616
rect 5592 6644 5598 6656
rect 5994 6644 6000 6656
rect 5592 6616 6000 6644
rect 5592 6604 5598 6616
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 8478 6604 8484 6656
rect 8536 6604 8542 6656
rect 10689 6647 10747 6653
rect 10689 6613 10701 6647
rect 10735 6644 10747 6647
rect 11238 6644 11244 6656
rect 10735 6616 11244 6644
rect 10735 6613 10747 6616
rect 10689 6607 10747 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11532 6644 11560 6820
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11977 6851 12035 6857
rect 11977 6848 11989 6851
rect 11664 6820 11989 6848
rect 11664 6808 11670 6820
rect 11977 6817 11989 6820
rect 12023 6817 12035 6851
rect 11977 6811 12035 6817
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 12124 6820 12173 6848
rect 12124 6808 12130 6820
rect 12161 6817 12173 6820
rect 12207 6848 12219 6851
rect 12250 6848 12256 6860
rect 12207 6820 12256 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12406 6848 12434 6888
rect 13188 6888 13492 6916
rect 12618 6848 12624 6860
rect 12406 6820 12624 6848
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 12802 6808 12808 6860
rect 12860 6808 12866 6860
rect 11609 6715 11667 6721
rect 11609 6681 11621 6715
rect 11655 6712 11667 6715
rect 13188 6712 13216 6888
rect 13262 6808 13268 6860
rect 13320 6808 13326 6860
rect 13464 6857 13492 6888
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13814 6848 13820 6860
rect 13495 6820 13820 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 15654 6848 15660 6860
rect 15243 6820 15660 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16301 6851 16359 6857
rect 16301 6848 16313 6851
rect 15988 6820 16313 6848
rect 15988 6808 15994 6820
rect 16301 6817 16313 6820
rect 16347 6817 16359 6851
rect 16301 6811 16359 6817
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16448 6820 16497 6848
rect 16448 6808 16454 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 16485 6811 16543 6817
rect 15378 6740 15384 6792
rect 15436 6740 15442 6792
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 15562 6740 15568 6792
rect 15620 6780 15626 6792
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 15620 6752 16129 6780
rect 15620 6740 15626 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 11655 6684 13216 6712
rect 11655 6681 11667 6684
rect 11609 6675 11667 6681
rect 11882 6644 11888 6656
rect 11532 6616 11888 6644
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 13446 6604 13452 6656
rect 13504 6604 13510 6656
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14700 6616 15025 6644
rect 14700 6604 14706 6616
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 15013 6607 15071 6613
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3660 6412 3985 6440
rect 3660 6400 3666 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 5442 6440 5448 6452
rect 3973 6403 4031 6409
rect 4540 6412 5448 6440
rect 3786 6264 3792 6316
rect 3844 6304 3850 6316
rect 4540 6313 4568 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5736 6412 6009 6440
rect 5258 6332 5264 6384
rect 5316 6372 5322 6384
rect 5736 6372 5764 6412
rect 5997 6409 6009 6412
rect 6043 6440 6055 6443
rect 7098 6440 7104 6452
rect 6043 6412 7104 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 8202 6400 8208 6452
rect 8260 6440 8266 6452
rect 8938 6440 8944 6452
rect 8260 6412 8944 6440
rect 8260 6400 8266 6412
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 11606 6400 11612 6452
rect 11664 6400 11670 6452
rect 11793 6443 11851 6449
rect 11793 6409 11805 6443
rect 11839 6440 11851 6443
rect 15562 6440 15568 6452
rect 11839 6412 15568 6440
rect 11839 6409 11851 6412
rect 11793 6403 11851 6409
rect 8294 6372 8300 6384
rect 5316 6344 5764 6372
rect 5828 6344 8300 6372
rect 5316 6332 5322 6344
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 3844 6276 4537 6304
rect 3844 6264 3850 6276
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 5718 6304 5724 6316
rect 4525 6267 4583 6273
rect 5184 6276 5724 6304
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 4893 6239 4951 6245
rect 4893 6236 4905 6239
rect 4856 6208 4905 6236
rect 4856 6196 4862 6208
rect 4893 6205 4905 6208
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 5074 6196 5080 6248
rect 5132 6196 5138 6248
rect 5184 6245 5212 6276
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5350 6236 5356 6248
rect 5307 6208 5356 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5828 6236 5856 6344
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6730 6304 6736 6316
rect 5960 6276 6736 6304
rect 5960 6264 5966 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 5500 6208 5856 6236
rect 5500 6196 5506 6208
rect 5994 6196 6000 6248
rect 6052 6196 6058 6248
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 7432 6208 7481 6236
rect 7432 6196 7438 6208
rect 7469 6205 7481 6208
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 7834 6236 7840 6248
rect 7791 6208 7840 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 7926 6196 7932 6248
rect 7984 6196 7990 6248
rect 8036 6245 8064 6344
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 11422 6332 11428 6384
rect 11480 6372 11486 6384
rect 11808 6372 11836 6403
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 16298 6400 16304 6452
rect 16356 6400 16362 6452
rect 11480 6344 11836 6372
rect 11480 6332 11486 6344
rect 12066 6332 12072 6384
rect 12124 6372 12130 6384
rect 12124 6344 13768 6372
rect 12124 6332 12130 6344
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8536 6276 10364 6304
rect 8536 6264 8542 6276
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 9674 6236 9680 6248
rect 8435 6208 9680 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10336 6236 10364 6276
rect 13170 6264 13176 6316
rect 13228 6304 13234 6316
rect 13740 6304 13768 6344
rect 14642 6332 14648 6384
rect 14700 6332 14706 6384
rect 15580 6372 15608 6400
rect 15580 6344 17080 6372
rect 15565 6307 15623 6313
rect 13228 6276 13676 6304
rect 13740 6276 14872 6304
rect 13228 6264 13234 6276
rect 10485 6239 10543 6245
rect 10485 6236 10497 6239
rect 10336 6208 10497 6236
rect 10229 6199 10287 6205
rect 10485 6205 10497 6208
rect 10531 6205 10543 6239
rect 10485 6199 10543 6205
rect 11701 6239 11759 6245
rect 11701 6205 11713 6239
rect 11747 6236 11759 6239
rect 11790 6236 11796 6248
rect 11747 6208 11796 6236
rect 11747 6205 11759 6208
rect 11701 6199 11759 6205
rect 4341 6171 4399 6177
rect 4341 6137 4353 6171
rect 4387 6168 4399 6171
rect 6178 6168 6184 6180
rect 4387 6140 6184 6168
rect 4387 6137 4399 6140
rect 4341 6131 4399 6137
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 8202 6168 8208 6180
rect 6288 6140 8208 6168
rect 4433 6103 4491 6109
rect 4433 6069 4445 6103
rect 4479 6100 4491 6103
rect 5534 6100 5540 6112
rect 4479 6072 5540 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 5534 6060 5540 6072
rect 5592 6060 5598 6112
rect 5626 6060 5632 6112
rect 5684 6060 5690 6112
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 6288 6100 6316 6140
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 10244 6168 10272 6199
rect 11790 6196 11796 6208
rect 11848 6196 11854 6248
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 9692 6140 10272 6168
rect 5868 6072 6316 6100
rect 5868 6060 5874 6072
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 8076 6072 8125 6100
rect 8076 6060 8082 6072
rect 8113 6069 8125 6072
rect 8159 6100 8171 6103
rect 8478 6100 8484 6112
rect 8159 6072 8484 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8478 6060 8484 6072
rect 8536 6060 8542 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 9692 6109 9720 6140
rect 11238 6128 11244 6180
rect 11296 6168 11302 6180
rect 13188 6168 13216 6264
rect 13538 6196 13544 6248
rect 13596 6196 13602 6248
rect 13648 6236 13676 6276
rect 13725 6239 13783 6245
rect 13725 6236 13737 6239
rect 13648 6208 13737 6236
rect 13725 6205 13737 6208
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 11296 6140 13216 6168
rect 13740 6168 13768 6199
rect 13814 6196 13820 6248
rect 13872 6196 13878 6248
rect 13906 6196 13912 6248
rect 13964 6196 13970 6248
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 14844 6245 14872 6276
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 15930 6304 15936 6316
rect 15611 6276 15936 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16448 6276 16589 6304
rect 16448 6264 16454 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 14332 6208 14565 6236
rect 14332 6196 14338 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 14737 6239 14795 6245
rect 14737 6205 14749 6239
rect 14783 6205 14795 6239
rect 14737 6199 14795 6205
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6205 14887 6239
rect 14829 6199 14887 6205
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15470 6236 15476 6248
rect 15243 6208 15476 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 14752 6168 14780 6199
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6205 15899 6239
rect 15841 6199 15899 6205
rect 15010 6168 15016 6180
rect 13740 6140 14688 6168
rect 14752 6140 15016 6168
rect 11296 6128 11302 6140
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9456 6072 9689 6100
rect 9456 6060 9462 6072
rect 9677 6069 9689 6072
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 13078 6100 13084 6112
rect 11848 6072 13084 6100
rect 11848 6060 11854 6072
rect 13078 6060 13084 6072
rect 13136 6100 13142 6112
rect 13814 6100 13820 6112
rect 13136 6072 13820 6100
rect 13136 6060 13142 6072
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14182 6060 14188 6112
rect 14240 6060 14246 6112
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 14332 6072 14381 6100
rect 14332 6060 14338 6072
rect 14369 6069 14381 6072
rect 14415 6069 14427 6103
rect 14660 6100 14688 6140
rect 15010 6128 15016 6140
rect 15068 6128 15074 6180
rect 15286 6128 15292 6180
rect 15344 6168 15350 6180
rect 15381 6171 15439 6177
rect 15381 6168 15393 6171
rect 15344 6140 15393 6168
rect 15344 6128 15350 6140
rect 15381 6137 15393 6140
rect 15427 6137 15439 6171
rect 15856 6168 15884 6199
rect 16022 6196 16028 6248
rect 16080 6196 16086 6248
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 17052 6245 17080 6344
rect 16485 6239 16543 6245
rect 16485 6205 16497 6239
rect 16531 6205 16543 6239
rect 16485 6199 16543 6205
rect 17037 6239 17095 6245
rect 17037 6205 17049 6239
rect 17083 6205 17095 6239
rect 17037 6199 17095 6205
rect 16500 6168 16528 6199
rect 16574 6168 16580 6180
rect 15856 6140 16580 6168
rect 15381 6131 15439 6137
rect 16574 6128 16580 6140
rect 16632 6128 16638 6180
rect 17218 6128 17224 6180
rect 17276 6128 17282 6180
rect 15194 6100 15200 6112
rect 14660 6072 15200 6100
rect 14369 6063 14427 6069
rect 15194 6060 15200 6072
rect 15252 6100 15258 6112
rect 16022 6100 16028 6112
rect 15252 6072 16028 6100
rect 15252 6060 15258 6072
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16945 6103 17003 6109
rect 16945 6100 16957 6103
rect 16448 6072 16957 6100
rect 16448 6060 16454 6072
rect 16945 6069 16957 6072
rect 16991 6100 17003 6103
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 16991 6072 17417 6100
rect 16991 6069 17003 6072
rect 16945 6063 17003 6069
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 5626 5896 5632 5908
rect 4632 5868 5632 5896
rect 3136 5763 3194 5769
rect 3136 5729 3148 5763
rect 3182 5760 3194 5763
rect 4062 5760 4068 5772
rect 3182 5732 4068 5760
rect 3182 5729 3194 5732
rect 3136 5723 3194 5729
rect 4062 5720 4068 5732
rect 4120 5760 4126 5772
rect 4632 5769 4660 5868
rect 5626 5856 5632 5868
rect 5684 5896 5690 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 5684 5868 6929 5896
rect 5684 5856 5690 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 7009 5899 7067 5905
rect 7009 5865 7021 5899
rect 7055 5896 7067 5899
rect 7055 5868 7604 5896
rect 7055 5865 7067 5868
rect 7009 5859 7067 5865
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 4847 5800 5212 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 4120 5732 4537 5760
rect 4120 5720 4126 5732
rect 4525 5729 4537 5732
rect 4571 5729 4583 5763
rect 4525 5723 4583 5729
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5729 4675 5763
rect 4617 5723 4675 5729
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 2884 5556 2912 5655
rect 4540 5624 4568 5723
rect 4890 5720 4896 5772
rect 4948 5720 4954 5772
rect 5074 5720 5080 5772
rect 5132 5720 5138 5772
rect 5184 5769 5212 5800
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 5592 5800 6101 5828
rect 5592 5788 5598 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 6181 5831 6239 5837
rect 6181 5797 6193 5831
rect 6227 5828 6239 5831
rect 7469 5831 7527 5837
rect 7469 5828 7481 5831
rect 6227 5800 7481 5828
rect 6227 5797 6239 5800
rect 6181 5791 6239 5797
rect 7469 5797 7481 5800
rect 7515 5797 7527 5831
rect 7469 5791 7527 5797
rect 7576 5772 7604 5868
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 9732 5868 11008 5896
rect 9732 5856 9738 5868
rect 10980 5837 11008 5868
rect 12526 5856 12532 5908
rect 12584 5896 12590 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12584 5868 12817 5896
rect 12584 5856 12590 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 14090 5896 14096 5908
rect 12805 5859 12863 5865
rect 13096 5868 14096 5896
rect 10965 5831 11023 5837
rect 10965 5797 10977 5831
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 13096 5772 13124 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 15010 5856 15016 5908
rect 15068 5856 15074 5908
rect 14274 5828 14280 5840
rect 13372 5800 14280 5828
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 5442 5720 5448 5772
rect 5500 5720 5506 5772
rect 5810 5720 5816 5772
rect 5868 5720 5874 5772
rect 5994 5769 6000 5772
rect 5961 5763 6000 5769
rect 5961 5729 5973 5763
rect 5961 5723 6000 5729
rect 5994 5720 6000 5723
rect 6052 5720 6058 5772
rect 6319 5763 6377 5769
rect 6319 5729 6331 5763
rect 6365 5760 6377 5763
rect 6365 5732 6776 5760
rect 6365 5729 6377 5732
rect 6319 5723 6377 5729
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 4982 5692 4988 5704
rect 4847 5664 4988 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 6178 5692 6184 5704
rect 5307 5664 6184 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 6748 5692 6776 5732
rect 6822 5720 6828 5772
rect 6880 5720 6886 5772
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7248 5732 7297 5760
rect 7248 5720 7254 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7374 5720 7380 5772
rect 7432 5720 7438 5772
rect 7558 5720 7564 5772
rect 7616 5720 7622 5772
rect 9306 5720 9312 5772
rect 9364 5720 9370 5772
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 9657 5763 9715 5769
rect 9657 5760 9669 5763
rect 9548 5732 9669 5760
rect 9548 5720 9554 5732
rect 9657 5729 9669 5732
rect 9703 5729 9715 5763
rect 9657 5723 9715 5729
rect 12986 5720 12992 5772
rect 13044 5720 13050 5772
rect 13078 5720 13084 5772
rect 13136 5720 13142 5772
rect 13170 5720 13176 5772
rect 13228 5720 13234 5772
rect 13372 5769 13400 5800
rect 14274 5788 14280 5800
rect 14332 5788 14338 5840
rect 14936 5828 14964 5856
rect 16853 5831 16911 5837
rect 16853 5828 16865 5831
rect 14936 5800 16252 5828
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 13446 5720 13452 5772
rect 13504 5760 13510 5772
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 13504 5732 13829 5760
rect 13504 5720 13510 5732
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 13998 5720 14004 5772
rect 14056 5720 14062 5772
rect 14185 5763 14243 5769
rect 14185 5729 14197 5763
rect 14231 5729 14243 5763
rect 14185 5723 14243 5729
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 14458 5760 14464 5772
rect 14415 5732 14464 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 7834 5692 7840 5704
rect 6748 5664 7840 5692
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8570 5692 8576 5704
rect 8352 5664 8576 5692
rect 8352 5652 8358 5664
rect 8570 5652 8576 5664
rect 8628 5692 8634 5704
rect 9398 5692 9404 5704
rect 8628 5664 9404 5692
rect 8628 5652 8634 5664
rect 9398 5652 9404 5664
rect 9456 5652 9462 5704
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 14016 5692 14044 5720
rect 13320 5664 14044 5692
rect 13320 5652 13326 5664
rect 7374 5624 7380 5636
rect 4540 5596 7380 5624
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 10781 5627 10839 5633
rect 10781 5593 10793 5627
rect 10827 5624 10839 5627
rect 11882 5624 11888 5636
rect 10827 5596 11888 5624
rect 10827 5593 10839 5596
rect 10781 5587 10839 5593
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 14200 5624 14228 5723
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 14921 5763 14979 5769
rect 14921 5729 14933 5763
rect 14967 5760 14979 5763
rect 15010 5760 15016 5772
rect 14967 5732 15016 5760
rect 14967 5729 14979 5732
rect 14921 5723 14979 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15105 5763 15163 5769
rect 15105 5729 15117 5763
rect 15151 5760 15163 5763
rect 15654 5760 15660 5772
rect 15151 5732 15660 5760
rect 15151 5729 15163 5732
rect 15105 5723 15163 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 16224 5769 16252 5800
rect 16592 5800 16865 5828
rect 16592 5772 16620 5800
rect 16853 5797 16865 5800
rect 16899 5797 16911 5831
rect 16853 5791 16911 5797
rect 16117 5763 16175 5769
rect 16117 5760 16129 5763
rect 16080 5732 16129 5760
rect 16080 5720 16086 5732
rect 16117 5729 16129 5732
rect 16163 5729 16175 5763
rect 16117 5723 16175 5729
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5729 16267 5763
rect 16209 5723 16267 5729
rect 16390 5720 16396 5772
rect 16448 5720 16454 5772
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 16574 5760 16580 5772
rect 16531 5732 16580 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16574 5720 16580 5732
rect 16632 5720 16638 5772
rect 16761 5763 16819 5769
rect 16761 5729 16773 5763
rect 16807 5729 16819 5763
rect 16761 5723 16819 5729
rect 16945 5763 17003 5769
rect 16945 5729 16957 5763
rect 16991 5760 17003 5763
rect 17218 5760 17224 5772
rect 16991 5732 17224 5760
rect 16991 5729 17003 5732
rect 16945 5723 17003 5729
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5692 14335 5695
rect 15470 5692 15476 5704
rect 14323 5664 15476 5692
rect 14323 5661 14335 5664
rect 14277 5655 14335 5661
rect 15470 5652 15476 5664
rect 15528 5692 15534 5704
rect 16776 5692 16804 5723
rect 15528 5664 16804 5692
rect 15528 5652 15534 5664
rect 13872 5596 14228 5624
rect 13872 5584 13878 5596
rect 15010 5584 15016 5636
rect 15068 5624 15074 5636
rect 15562 5624 15568 5636
rect 15068 5596 15568 5624
rect 15068 5584 15074 5596
rect 15562 5584 15568 5596
rect 15620 5584 15626 5636
rect 16206 5584 16212 5636
rect 16264 5624 16270 5636
rect 16960 5624 16988 5723
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 16264 5596 16988 5624
rect 16264 5584 16270 5596
rect 3970 5556 3976 5568
rect 2884 5528 3976 5556
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5534 5556 5540 5568
rect 4948 5528 5540 5556
rect 4948 5516 4954 5528
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5629 5559 5687 5565
rect 5629 5525 5641 5559
rect 5675 5556 5687 5559
rect 5810 5556 5816 5568
rect 5675 5528 5816 5556
rect 5675 5525 5687 5528
rect 5629 5519 5687 5525
rect 5810 5516 5816 5528
rect 5868 5516 5874 5568
rect 6454 5516 6460 5568
rect 6512 5516 6518 5568
rect 6546 5516 6552 5568
rect 6604 5516 6610 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7193 5559 7251 5565
rect 7193 5556 7205 5559
rect 7156 5528 7205 5556
rect 7156 5516 7162 5528
rect 7193 5525 7205 5528
rect 7239 5556 7251 5559
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 7239 5528 9229 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 9217 5525 9229 5528
rect 9263 5556 9275 5559
rect 9398 5556 9404 5568
rect 9263 5528 9404 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11422 5516 11428 5568
rect 11480 5556 11486 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 11480 5528 12265 5556
rect 11480 5516 11486 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14642 5556 14648 5568
rect 13955 5528 14648 5556
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 14976 5528 16681 5556
rect 14976 5516 14982 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 16669 5519 16727 5525
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6454 5352 6460 5364
rect 6227 5324 6460 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6696 5324 8064 5352
rect 6696 5312 6702 5324
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 7745 5287 7803 5293
rect 7745 5284 7757 5287
rect 5132 5256 7757 5284
rect 5132 5244 5138 5256
rect 6273 5219 6331 5225
rect 6273 5185 6285 5219
rect 6319 5216 6331 5219
rect 6546 5216 6552 5228
rect 6319 5188 6552 5216
rect 6319 5185 6331 5188
rect 6273 5179 6331 5185
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 5810 5151 5868 5157
rect 5810 5117 5822 5151
rect 5856 5148 5868 5151
rect 6914 5148 6920 5160
rect 5856 5120 6920 5148
rect 5856 5117 5868 5120
rect 5810 5111 5868 5117
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 7668 5157 7696 5256
rect 7745 5253 7757 5256
rect 7791 5253 7803 5287
rect 7745 5247 7803 5253
rect 8036 5284 8064 5324
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11974 5352 11980 5364
rect 11112 5324 11980 5352
rect 11112 5312 11118 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12894 5312 12900 5364
rect 12952 5312 12958 5364
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 13228 5324 14289 5352
rect 13228 5312 13234 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 15470 5312 15476 5364
rect 15528 5312 15534 5364
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 16301 5355 16359 5361
rect 16301 5352 16313 5355
rect 16080 5324 16313 5352
rect 16080 5312 16086 5324
rect 16301 5321 16313 5324
rect 16347 5321 16359 5355
rect 16301 5315 16359 5321
rect 8478 5284 8484 5296
rect 8036 5256 8484 5284
rect 7469 5151 7527 5157
rect 7469 5148 7481 5151
rect 7340 5120 7481 5148
rect 7340 5108 7346 5120
rect 7469 5117 7481 5120
rect 7515 5117 7527 5151
rect 7469 5111 7527 5117
rect 7653 5151 7711 5157
rect 7653 5117 7665 5151
rect 7699 5148 7711 5151
rect 7742 5148 7748 5160
rect 7699 5120 7748 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8036 5148 8064 5256
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 8570 5244 8576 5296
rect 8628 5284 8634 5296
rect 11146 5284 11152 5296
rect 8628 5256 11152 5284
rect 8628 5244 8634 5256
rect 11146 5244 11152 5256
rect 11204 5284 11210 5296
rect 11425 5287 11483 5293
rect 11425 5284 11437 5287
rect 11204 5256 11437 5284
rect 11204 5244 11210 5256
rect 11425 5253 11437 5256
rect 11471 5253 11483 5287
rect 11425 5247 11483 5253
rect 12802 5244 12808 5296
rect 12860 5284 12866 5296
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 12860 5256 14504 5284
rect 12860 5244 12866 5256
rect 8662 5216 8668 5228
rect 8220 5188 8668 5216
rect 8220 5157 8248 5188
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10928 5188 11376 5216
rect 10928 5176 10934 5188
rect 7975 5120 8064 5148
rect 8205 5151 8263 5157
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 8205 5117 8217 5151
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 8536 5120 8585 5148
rect 8536 5108 8542 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8757 5151 8815 5157
rect 8757 5117 8769 5151
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 8938 5148 8944 5160
rect 8895 5120 8944 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6638 5080 6644 5092
rect 6052 5052 6644 5080
rect 6052 5040 6058 5052
rect 6638 5040 6644 5052
rect 6696 5040 6702 5092
rect 7561 5083 7619 5089
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 8113 5083 8171 5089
rect 7607 5052 7880 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 5810 4972 5816 5024
rect 5868 4972 5874 5024
rect 7852 5012 7880 5052
rect 8113 5049 8125 5083
rect 8159 5080 8171 5083
rect 8772 5080 8800 5111
rect 8938 5108 8944 5120
rect 8996 5108 9002 5160
rect 11238 5108 11244 5160
rect 11296 5108 11302 5160
rect 11348 5157 11376 5188
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12621 5219 12679 5225
rect 12124 5188 12572 5216
rect 12124 5176 12130 5188
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5117 11391 5151
rect 11333 5111 11391 5117
rect 12434 5108 12440 5160
rect 12492 5108 12498 5160
rect 12544 5157 12572 5188
rect 12621 5185 12633 5219
rect 12667 5216 12679 5219
rect 14366 5216 14372 5228
rect 12667 5188 14372 5216
rect 12667 5185 12679 5188
rect 12621 5179 12679 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 12529 5151 12587 5157
rect 12529 5117 12541 5151
rect 12575 5117 12587 5151
rect 12529 5111 12587 5117
rect 11054 5080 11060 5092
rect 8159 5052 8524 5080
rect 8159 5049 8171 5052
rect 8113 5043 8171 5049
rect 7926 5012 7932 5024
rect 7852 4984 7932 5012
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8076 4984 8401 5012
rect 8076 4972 8082 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8496 5012 8524 5052
rect 8772 5052 11060 5080
rect 8772 5012 8800 5052
rect 11054 5040 11060 5052
rect 11112 5040 11118 5092
rect 12544 5080 12572 5111
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5148 13047 5151
rect 13814 5148 13820 5160
rect 13035 5120 13820 5148
rect 13035 5117 13047 5120
rect 12989 5111 13047 5117
rect 13004 5080 13032 5111
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14182 5108 14188 5160
rect 14240 5108 14246 5160
rect 14476 5157 14504 5256
rect 14568 5256 16129 5284
rect 14568 5225 14596 5256
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 14918 5176 14924 5228
rect 14976 5176 14982 5228
rect 15378 5216 15384 5228
rect 15028 5188 15384 5216
rect 14461 5151 14519 5157
rect 14461 5117 14473 5151
rect 14507 5148 14519 5151
rect 15028 5148 15056 5188
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 14507 5120 15056 5148
rect 14507 5117 14519 5120
rect 14461 5111 14519 5117
rect 15194 5108 15200 5160
rect 15252 5108 15258 5160
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15565 5151 15623 5157
rect 15565 5148 15577 5151
rect 15528 5120 15577 5148
rect 15528 5108 15534 5120
rect 15565 5117 15577 5120
rect 15611 5148 15623 5151
rect 16206 5148 16212 5160
rect 15611 5120 16212 5148
rect 15611 5117 15623 5120
rect 15565 5111 15623 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 16298 5108 16304 5160
rect 16356 5108 16362 5160
rect 16482 5108 16488 5160
rect 16540 5108 16546 5160
rect 14829 5083 14887 5089
rect 14829 5080 14841 5083
rect 12544 5052 13032 5080
rect 14384 5052 14841 5080
rect 14384 5024 14412 5052
rect 14829 5049 14841 5052
rect 14875 5049 14887 5083
rect 14829 5043 14887 5049
rect 8496 4984 8800 5012
rect 8389 4975 8447 4981
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 12894 5012 12900 5024
rect 11572 4984 12900 5012
rect 11572 4972 11578 4984
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13078 4972 13084 5024
rect 13136 4972 13142 5024
rect 14090 4972 14096 5024
rect 14148 4972 14154 5024
rect 14366 4972 14372 5024
rect 14424 4972 14430 5024
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 14918 5012 14924 5024
rect 14700 4984 14924 5012
rect 14700 4972 14706 4984
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15010 4972 15016 5024
rect 15068 4972 15074 5024
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 6273 4811 6331 4817
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 6914 4808 6920 4820
rect 6319 4780 6920 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7834 4808 7840 4820
rect 7300 4780 7840 4808
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6362 4672 6368 4684
rect 6319 4644 6368 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6104 4604 6132 4635
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7300 4681 7328 4780
rect 7834 4768 7840 4780
rect 7892 4808 7898 4820
rect 7892 4780 8708 4808
rect 7892 4768 7898 4780
rect 7374 4700 7380 4752
rect 7432 4740 7438 4752
rect 7432 4712 7696 4740
rect 7432 4700 7438 4712
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 7208 4604 7236 4635
rect 7392 4604 7420 4700
rect 7561 4675 7619 4681
rect 7561 4641 7573 4675
rect 7607 4641 7619 4675
rect 7561 4635 7619 4641
rect 6104 4576 7420 4604
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 7377 4539 7435 4545
rect 7377 4505 7389 4539
rect 7423 4536 7435 4539
rect 7576 4536 7604 4635
rect 7668 4604 7696 4712
rect 8570 4700 8576 4752
rect 8628 4700 8634 4752
rect 7742 4632 7748 4684
rect 7800 4632 7806 4684
rect 7834 4632 7840 4684
rect 7892 4632 7898 4684
rect 7926 4632 7932 4684
rect 7984 4632 7990 4684
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4672 8079 4675
rect 8386 4672 8392 4684
rect 8067 4644 8392 4672
rect 8067 4641 8079 4644
rect 8021 4635 8079 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8481 4675 8539 4681
rect 8481 4641 8493 4675
rect 8527 4672 8539 4675
rect 8588 4672 8616 4700
rect 8680 4681 8708 4780
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 11057 4811 11115 4817
rect 11057 4808 11069 4811
rect 11020 4780 11069 4808
rect 11020 4768 11026 4780
rect 11057 4777 11069 4780
rect 11103 4808 11115 4811
rect 12342 4808 12348 4820
rect 11103 4780 12348 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12434 4768 12440 4820
rect 12492 4768 12498 4820
rect 12710 4768 12716 4820
rect 12768 4768 12774 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 14274 4808 14280 4820
rect 12952 4780 14280 4808
rect 12952 4768 12958 4780
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14516 4780 14841 4808
rect 14516 4768 14522 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 14829 4771 14887 4777
rect 13078 4740 13084 4752
rect 12360 4712 13084 4740
rect 8527 4644 8616 4672
rect 8665 4675 8723 4681
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 8665 4641 8677 4675
rect 8711 4641 8723 4675
rect 8665 4635 8723 4641
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 10928 4644 11253 4672
rect 10928 4632 10934 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 11241 4635 11299 4641
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4672 11483 4675
rect 11514 4672 11520 4684
rect 11471 4644 11520 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 7668 4576 8585 4604
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 11256 4604 11284 4635
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 11701 4675 11759 4681
rect 11701 4641 11713 4675
rect 11747 4641 11759 4675
rect 11701 4635 11759 4641
rect 11716 4604 11744 4635
rect 11974 4632 11980 4684
rect 12032 4672 12038 4684
rect 12253 4675 12311 4681
rect 12253 4672 12265 4675
rect 12032 4644 12265 4672
rect 12032 4632 12038 4644
rect 12253 4641 12265 4644
rect 12299 4641 12311 4675
rect 12253 4635 12311 4641
rect 11256 4576 11744 4604
rect 12069 4607 12127 4613
rect 8573 4567 8631 4573
rect 12069 4573 12081 4607
rect 12115 4604 12127 4607
rect 12360 4604 12388 4712
rect 13078 4700 13084 4712
rect 13136 4700 13142 4752
rect 14292 4740 14320 4768
rect 14200 4712 14320 4740
rect 15105 4743 15163 4749
rect 12710 4632 12716 4684
rect 12768 4632 12774 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 14090 4672 14096 4684
rect 12943 4644 14096 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 14200 4681 14228 4712
rect 15105 4709 15117 4743
rect 15151 4740 15163 4743
rect 15657 4743 15715 4749
rect 15657 4740 15669 4743
rect 15151 4712 15669 4740
rect 15151 4709 15163 4712
rect 15105 4703 15163 4709
rect 15657 4709 15669 4712
rect 15703 4709 15715 4743
rect 15657 4703 15715 4709
rect 14185 4675 14243 4681
rect 14185 4641 14197 4675
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14369 4675 14427 4681
rect 14369 4672 14381 4675
rect 14332 4644 14381 4672
rect 14332 4632 14338 4644
rect 14369 4641 14381 4644
rect 14415 4641 14427 4675
rect 14369 4635 14427 4641
rect 14550 4632 14556 4684
rect 14608 4632 14614 4684
rect 14734 4632 14740 4684
rect 14792 4632 14798 4684
rect 14918 4632 14924 4684
rect 14976 4681 14982 4684
rect 14976 4675 15025 4681
rect 14976 4641 14979 4675
rect 15013 4641 15025 4675
rect 14976 4635 15025 4641
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 15380 4675 15438 4681
rect 15380 4641 15392 4675
rect 15426 4641 15438 4675
rect 15380 4635 15438 4641
rect 14976 4632 14982 4635
rect 12115 4576 12388 4604
rect 12115 4573 12127 4576
rect 12069 4567 12127 4573
rect 12434 4564 12440 4616
rect 12492 4604 12498 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12492 4576 12817 4604
rect 12492 4564 12498 4576
rect 12805 4573 12817 4576
rect 12851 4604 12863 4607
rect 12851 4576 13032 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 11517 4539 11575 4545
rect 7423 4508 8432 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8404 4480 8432 4508
rect 11517 4505 11529 4539
rect 11563 4536 11575 4539
rect 12710 4536 12716 4548
rect 11563 4508 12716 4536
rect 11563 4505 11575 4508
rect 11517 4499 11575 4505
rect 12710 4496 12716 4508
rect 12768 4496 12774 4548
rect 8202 4428 8208 4480
rect 8260 4428 8266 4480
rect 8386 4428 8392 4480
rect 8444 4428 8450 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8849 4471 8907 4477
rect 8849 4468 8861 4471
rect 8720 4440 8861 4468
rect 8720 4428 8726 4440
rect 8849 4437 8861 4440
rect 8895 4437 8907 4471
rect 8849 4431 8907 4437
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 12894 4468 12900 4480
rect 11931 4440 12900 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13004 4468 13032 4576
rect 13170 4564 13176 4616
rect 13228 4564 13234 4616
rect 13998 4564 14004 4616
rect 14056 4564 14062 4616
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14568 4604 14596 4632
rect 15212 4604 15240 4635
rect 14568 4576 15240 4604
rect 15395 4604 15423 4635
rect 15470 4632 15476 4684
rect 15528 4632 15534 4684
rect 15562 4632 15568 4684
rect 15620 4632 15626 4684
rect 15749 4675 15807 4681
rect 15749 4641 15761 4675
rect 15795 4672 15807 4675
rect 16114 4672 16120 4684
rect 15795 4644 16120 4672
rect 15795 4641 15807 4644
rect 15749 4635 15807 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 15580 4604 15608 4632
rect 15395 4576 15608 4604
rect 13081 4539 13139 4545
rect 13081 4505 13093 4539
rect 13127 4536 13139 4539
rect 13538 4536 13544 4548
rect 13127 4508 13544 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 13538 4496 13544 4508
rect 13596 4496 13602 4548
rect 13814 4496 13820 4548
rect 13872 4536 13878 4548
rect 14734 4536 14740 4548
rect 13872 4508 14740 4536
rect 13872 4496 13878 4508
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 15395 4468 15423 4576
rect 13004 4440 15423 4468
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 8662 4224 8668 4276
rect 8720 4224 8726 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12253 4267 12311 4273
rect 12253 4264 12265 4267
rect 12032 4236 12265 4264
rect 12032 4224 12038 4236
rect 12253 4233 12265 4236
rect 12299 4233 12311 4267
rect 12253 4227 12311 4233
rect 12894 4224 12900 4276
rect 12952 4264 12958 4276
rect 13722 4264 13728 4276
rect 12952 4236 13728 4264
rect 12952 4224 12958 4236
rect 13722 4224 13728 4236
rect 13780 4264 13786 4276
rect 14001 4267 14059 4273
rect 13780 4236 13952 4264
rect 13780 4224 13786 4236
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 8938 4196 8944 4208
rect 7432 4168 8944 4196
rect 7432 4156 7438 4168
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 13814 4196 13820 4208
rect 13096 4168 13820 4196
rect 3970 4020 3976 4072
rect 4028 4060 4034 4072
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 4028 4032 5825 4060
rect 4028 4020 4034 4032
rect 5813 4029 5825 4032
rect 5859 4060 5871 4063
rect 8294 4060 8300 4072
rect 5859 4032 8300 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8386 4020 8392 4072
rect 8444 4020 8450 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 9355 4032 10885 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 10873 4029 10885 4032
rect 10919 4060 10931 4063
rect 11422 4060 11428 4072
rect 10919 4032 11428 4060
rect 10919 4029 10931 4032
rect 10873 4023 10931 4029
rect 11422 4020 11428 4032
rect 11480 4020 11486 4072
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4029 12587 4063
rect 12529 4023 12587 4029
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 6058 3995 6116 4001
rect 6058 3992 6070 3995
rect 5684 3964 6070 3992
rect 5684 3952 5690 3964
rect 6058 3961 6070 3964
rect 6104 3961 6116 3995
rect 6058 3955 6116 3961
rect 8938 3952 8944 4004
rect 8996 3992 9002 4004
rect 11146 4001 11152 4004
rect 9554 3995 9612 4001
rect 9554 3992 9566 3995
rect 8996 3964 9566 3992
rect 8996 3952 9002 3964
rect 9554 3961 9566 3964
rect 9600 3961 9612 3995
rect 9554 3955 9612 3961
rect 11140 3955 11152 4001
rect 11146 3952 11152 3955
rect 11204 3952 11210 4004
rect 11330 3952 11336 4004
rect 11388 3992 11394 4004
rect 12345 3995 12403 4001
rect 12345 3992 12357 3995
rect 11388 3964 12357 3992
rect 11388 3952 11394 3964
rect 12345 3961 12357 3964
rect 12391 3961 12403 3995
rect 12544 3992 12572 4023
rect 12802 4020 12808 4072
rect 12860 4020 12866 4072
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13096 4060 13124 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 13924 4196 13952 4236
rect 14001 4233 14013 4267
rect 14047 4264 14059 4267
rect 14458 4264 14464 4276
rect 14047 4236 14464 4264
rect 14047 4233 14059 4236
rect 14001 4227 14059 4233
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 16298 4196 16304 4208
rect 13924 4168 16304 4196
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13228 4100 13645 4128
rect 13228 4088 13234 4100
rect 13633 4097 13645 4100
rect 13679 4097 13691 4131
rect 14918 4128 14924 4140
rect 13633 4091 13691 4097
rect 14476 4100 14924 4128
rect 13035 4032 13124 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 13722 4020 13728 4072
rect 13780 4020 13786 4072
rect 14476 4069 14504 4100
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 14645 4063 14703 4069
rect 14645 4029 14657 4063
rect 14691 4060 14703 4063
rect 15010 4060 15016 4072
rect 14691 4032 15016 4060
rect 14691 4029 14703 4032
rect 14645 4023 14703 4029
rect 15010 4020 15016 4032
rect 15068 4020 15074 4072
rect 13998 3992 14004 4004
rect 12544 3964 14004 3992
rect 12345 3955 12403 3961
rect 13998 3952 14004 3964
rect 14056 3952 14062 4004
rect 7190 3884 7196 3936
rect 7248 3884 7254 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9674 3924 9680 3936
rect 8895 3896 9680 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10689 3927 10747 3933
rect 10689 3893 10701 3927
rect 10735 3924 10747 3927
rect 11514 3924 11520 3936
rect 10735 3896 11520 3924
rect 10735 3893 10747 3896
rect 10689 3887 10747 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 9861 3723 9919 3729
rect 9861 3689 9873 3723
rect 9907 3720 9919 3723
rect 10870 3720 10876 3732
rect 9907 3692 10876 3720
rect 9907 3689 9919 3692
rect 9861 3683 9919 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 12345 3723 12403 3729
rect 12345 3689 12357 3723
rect 12391 3720 12403 3723
rect 12802 3720 12808 3732
rect 12391 3692 12808 3720
rect 12391 3689 12403 3692
rect 12345 3683 12403 3689
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 7190 3612 7196 3664
rect 7248 3652 7254 3664
rect 11054 3652 11060 3664
rect 7248 3624 10088 3652
rect 7248 3612 7254 3624
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 8352 3556 8493 3584
rect 8352 3544 8358 3556
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 8748 3587 8806 3593
rect 8748 3584 8760 3587
rect 8628 3556 8760 3584
rect 8628 3544 8634 3556
rect 8748 3553 8760 3556
rect 8794 3553 8806 3587
rect 8748 3547 8806 3553
rect 9674 3544 9680 3596
rect 9732 3584 9738 3596
rect 9953 3587 10011 3593
rect 9953 3584 9965 3587
rect 9732 3556 9965 3584
rect 9732 3544 9738 3556
rect 9953 3553 9965 3556
rect 9999 3553 10011 3587
rect 9953 3547 10011 3553
rect 10060 3380 10088 3624
rect 10980 3624 11060 3652
rect 10980 3593 11008 3624
rect 11054 3612 11060 3624
rect 11112 3652 11118 3664
rect 11422 3652 11428 3664
rect 11112 3624 11428 3652
rect 11112 3612 11118 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 10965 3587 11023 3593
rect 10965 3553 10977 3587
rect 11011 3553 11023 3587
rect 11221 3587 11279 3593
rect 11221 3584 11233 3587
rect 10965 3547 11023 3553
rect 11072 3556 11233 3584
rect 11072 3516 11100 3556
rect 11221 3553 11233 3556
rect 11267 3553 11279 3587
rect 11221 3547 11279 3553
rect 10152 3488 11100 3516
rect 10152 3457 10180 3488
rect 10137 3451 10195 3457
rect 10137 3417 10149 3451
rect 10183 3417 10195 3451
rect 10137 3411 10195 3417
rect 12986 3380 12992 3392
rect 10060 3352 12992 3380
rect 12986 3340 12992 3352
rect 13044 3340 13050 3392
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 3694 2864 3700 2916
rect 3752 2904 3758 2916
rect 3752 2876 12434 2904
rect 3752 2864 3758 2876
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 11790 2836 11796 2848
rect 6236 2808 11796 2836
rect 6236 2796 6242 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12406 2836 12434 2876
rect 12802 2836 12808 2848
rect 12406 2808 12808 2836
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8662 2632 8668 2644
rect 7791 2604 8668 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 12802 2592 12808 2644
rect 12860 2592 12866 2644
rect 8880 2567 8938 2573
rect 8880 2533 8892 2567
rect 8926 2564 8938 2567
rect 10226 2564 10232 2576
rect 8926 2536 10232 2564
rect 8926 2533 8938 2536
rect 8880 2527 8938 2533
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 13940 2567 13998 2573
rect 13940 2533 13952 2567
rect 13986 2564 13998 2567
rect 15102 2564 15108 2576
rect 13986 2536 15108 2564
rect 13986 2533 13998 2536
rect 13940 2527 13998 2533
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 11054 2428 11060 2440
rect 9171 2400 11060 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2428 14243 2431
rect 14274 2428 14280 2440
rect 14231 2400 14280 2428
rect 14231 2397 14243 2400
rect 14185 2391 14243 2397
rect 14274 2388 14280 2400
rect 14332 2388 14338 2440
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 10045 1887 10103 1893
rect 10045 1853 10057 1887
rect 10091 1884 10103 1887
rect 11054 1884 11060 1896
rect 10091 1856 11060 1884
rect 10091 1853 10103 1856
rect 10045 1847 10103 1853
rect 11054 1844 11060 1856
rect 11112 1844 11118 1896
rect 10312 1819 10370 1825
rect 10312 1785 10324 1819
rect 10358 1816 10370 1819
rect 10594 1816 10600 1828
rect 10358 1788 10600 1816
rect 10358 1785 10370 1788
rect 10312 1779 10370 1785
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 11425 1751 11483 1757
rect 11425 1748 11437 1751
rect 11204 1720 11437 1748
rect 11204 1708 11210 1720
rect 11425 1717 11437 1720
rect 11471 1717 11483 1751
rect 11425 1711 11483 1717
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 1210 1504 1216 1556
rect 1268 1544 1274 1556
rect 2593 1547 2651 1553
rect 2593 1544 2605 1547
rect 1268 1516 2605 1544
rect 1268 1504 1274 1516
rect 2593 1513 2605 1516
rect 2639 1513 2651 1547
rect 2593 1507 2651 1513
rect 11790 1504 11796 1556
rect 11848 1504 11854 1556
rect 13630 1504 13636 1556
rect 13688 1544 13694 1556
rect 14645 1547 14703 1553
rect 14645 1544 14657 1547
rect 13688 1516 14657 1544
rect 13688 1504 13694 1516
rect 14645 1513 14657 1516
rect 14691 1513 14703 1547
rect 14645 1507 14703 1513
rect 16666 1504 16672 1556
rect 16724 1544 16730 1556
rect 17865 1547 17923 1553
rect 16724 1516 16804 1544
rect 16724 1504 16730 1516
rect 11698 1436 11704 1488
rect 11756 1476 11762 1488
rect 12906 1479 12964 1485
rect 12906 1476 12918 1479
rect 11756 1448 12918 1476
rect 11756 1436 11762 1448
rect 12906 1445 12918 1448
rect 12952 1445 12964 1479
rect 12906 1439 12964 1445
rect 13078 1436 13084 1488
rect 13136 1476 13142 1488
rect 16776 1485 16804 1516
rect 17865 1513 17877 1547
rect 17911 1544 17923 1547
rect 18598 1544 18604 1556
rect 17911 1516 18604 1544
rect 17911 1513 17923 1516
rect 17865 1507 17923 1513
rect 18598 1504 18604 1516
rect 18656 1504 18662 1556
rect 13510 1479 13568 1485
rect 13510 1476 13522 1479
rect 13136 1448 13522 1476
rect 13136 1436 13142 1448
rect 13510 1445 13522 1448
rect 13556 1445 13568 1479
rect 13510 1439 13568 1445
rect 16752 1479 16810 1485
rect 16752 1445 16764 1479
rect 16798 1445 16810 1479
rect 16752 1439 16810 1445
rect 3717 1411 3775 1417
rect 3717 1408 3729 1411
rect 2976 1380 3729 1408
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1340 2283 1343
rect 2976 1340 3004 1380
rect 3717 1377 3729 1380
rect 3763 1408 3775 1411
rect 3878 1408 3884 1420
rect 3763 1380 3884 1408
rect 3763 1377 3775 1380
rect 3717 1371 3775 1377
rect 3878 1368 3884 1380
rect 3936 1368 3942 1420
rect 11054 1368 11060 1420
rect 11112 1408 11118 1420
rect 13814 1408 13820 1420
rect 11112 1380 13820 1408
rect 11112 1368 11118 1380
rect 2271 1312 3004 1340
rect 2271 1309 2283 1312
rect 2225 1303 2283 1309
rect 3970 1300 3976 1352
rect 4028 1300 4034 1352
rect 13280 1349 13308 1380
rect 13814 1368 13820 1380
rect 13872 1408 13878 1420
rect 14274 1408 14280 1420
rect 13872 1380 14280 1408
rect 13872 1368 13878 1380
rect 14274 1368 14280 1380
rect 14332 1368 14338 1420
rect 13173 1343 13231 1349
rect 13173 1309 13185 1343
rect 13219 1340 13231 1343
rect 13265 1343 13323 1349
rect 13265 1340 13277 1343
rect 13219 1312 13277 1340
rect 13219 1309 13231 1312
rect 13173 1303 13231 1309
rect 13265 1309 13277 1312
rect 13311 1309 13323 1343
rect 14292 1340 14320 1368
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 14292 1312 16497 1340
rect 13265 1303 13323 1309
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16485 1303 16543 1309
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 13814 1000 13820 1012
rect 13648 972 13820 1000
rect 13648 873 13676 972
rect 13814 960 13820 972
rect 13872 960 13878 1012
rect 13633 867 13691 873
rect 13633 833 13645 867
rect 13679 833 13691 867
rect 13633 827 13691 833
rect 13906 805 13912 808
rect 13900 759 13912 805
rect 13906 756 13912 759
rect 13964 756 13970 808
rect 15013 663 15071 669
rect 15013 629 15025 663
rect 15059 660 15071 663
rect 16114 660 16120 672
rect 15059 632 16120 660
rect 15059 629 15071 632
rect 15013 623 15071 629
rect 16114 620 16120 632
rect 16172 620 16178 672
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 10508 18912 10560 18964
rect 8392 18844 8444 18896
rect 848 18776 900 18828
rect 2504 18776 2556 18828
rect 4160 18776 4212 18828
rect 5816 18776 5868 18828
rect 6368 18819 6420 18828
rect 6368 18785 6377 18819
rect 6377 18785 6411 18819
rect 6411 18785 6420 18819
rect 6368 18776 6420 18785
rect 7472 18776 7524 18828
rect 9128 18776 9180 18828
rect 10784 18776 10836 18828
rect 12440 18776 12492 18828
rect 14096 18776 14148 18828
rect 15752 18776 15804 18828
rect 17408 18776 17460 18828
rect 10140 18640 10192 18692
rect 5908 18572 5960 18624
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 8024 18572 8076 18624
rect 10416 18640 10468 18692
rect 12532 18640 12584 18692
rect 10324 18572 10376 18624
rect 11980 18572 12032 18624
rect 12808 18572 12860 18624
rect 13544 18572 13596 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16672 18572 16724 18624
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 11888 18411 11940 18420
rect 7380 18232 7432 18284
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 9680 18300 9732 18352
rect 10784 18300 10836 18352
rect 4252 18096 4304 18148
rect 4712 18096 4764 18148
rect 5448 18096 5500 18148
rect 5632 18096 5684 18148
rect 6092 18139 6144 18148
rect 6092 18105 6126 18139
rect 6126 18105 6144 18139
rect 6092 18096 6144 18105
rect 6276 18096 6328 18148
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 12072 18164 12124 18216
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 8484 18096 8536 18148
rect 11060 18096 11112 18148
rect 12624 18096 12676 18148
rect 8208 18071 8260 18080
rect 8208 18037 8217 18071
rect 8217 18037 8251 18071
rect 8251 18037 8260 18071
rect 8208 18028 8260 18037
rect 9588 18028 9640 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 16580 18071 16632 18080
rect 16580 18037 16589 18071
rect 16589 18037 16623 18071
rect 16623 18037 16632 18071
rect 16580 18028 16632 18037
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 4252 17867 4304 17876
rect 4252 17833 4261 17867
rect 4261 17833 4295 17867
rect 4295 17833 4304 17867
rect 4252 17824 4304 17833
rect 6368 17824 6420 17876
rect 7380 17867 7432 17876
rect 4804 17756 4856 17808
rect 7380 17833 7407 17867
rect 7407 17833 7432 17867
rect 7380 17824 7432 17833
rect 8484 17824 8536 17876
rect 5448 17620 5500 17672
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 4712 17527 4764 17536
rect 4712 17493 4721 17527
rect 4721 17493 4755 17527
rect 4755 17493 4764 17527
rect 4712 17484 4764 17493
rect 5632 17552 5684 17604
rect 7840 17756 7892 17808
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 9680 17688 9732 17740
rect 10600 17824 10652 17876
rect 11060 17824 11112 17876
rect 12624 17867 12676 17876
rect 12624 17833 12633 17867
rect 12633 17833 12667 17867
rect 12667 17833 12676 17867
rect 12624 17824 12676 17833
rect 10324 17620 10376 17672
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 12808 17731 12860 17740
rect 12808 17697 12817 17731
rect 12817 17697 12851 17731
rect 12851 17697 12860 17731
rect 12808 17688 12860 17697
rect 12900 17731 12952 17740
rect 12900 17697 12909 17731
rect 12909 17697 12943 17731
rect 12943 17697 12952 17731
rect 12900 17688 12952 17697
rect 10784 17620 10836 17672
rect 5540 17484 5592 17536
rect 11060 17552 11112 17604
rect 15108 17620 15160 17672
rect 7380 17527 7432 17536
rect 7380 17493 7389 17527
rect 7389 17493 7423 17527
rect 7423 17493 7432 17527
rect 7380 17484 7432 17493
rect 9220 17527 9272 17536
rect 9220 17493 9229 17527
rect 9229 17493 9263 17527
rect 9263 17493 9272 17527
rect 9220 17484 9272 17493
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 5724 17280 5776 17332
rect 8116 17323 8168 17332
rect 8116 17289 8125 17323
rect 8125 17289 8159 17323
rect 8159 17289 8168 17323
rect 8116 17280 8168 17289
rect 12348 17280 12400 17332
rect 7012 17212 7064 17264
rect 7840 17212 7892 17264
rect 4804 17076 4856 17128
rect 8116 17076 8168 17128
rect 5448 17008 5500 17060
rect 7380 17008 7432 17060
rect 9680 17212 9732 17264
rect 10232 17144 10284 17196
rect 10600 17144 10652 17196
rect 11612 17144 11664 17196
rect 12900 17212 12952 17264
rect 10968 17076 11020 17128
rect 12256 17144 12308 17196
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 4988 16983 5040 16992
rect 4988 16949 4997 16983
rect 4997 16949 5031 16983
rect 5031 16949 5040 16983
rect 4988 16940 5040 16949
rect 5632 16940 5684 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 11060 17008 11112 17060
rect 9128 16940 9180 16992
rect 10416 16940 10468 16992
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 16580 17076 16632 17128
rect 13544 17008 13596 17060
rect 12624 16940 12676 16992
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 7380 16736 7432 16788
rect 2320 16600 2372 16652
rect 4344 16600 4396 16652
rect 5540 16643 5592 16652
rect 5540 16609 5549 16643
rect 5549 16609 5583 16643
rect 5583 16609 5592 16643
rect 5540 16600 5592 16609
rect 6276 16643 6328 16652
rect 6276 16609 6285 16643
rect 6285 16609 6319 16643
rect 6319 16609 6328 16643
rect 6276 16600 6328 16609
rect 6552 16643 6604 16652
rect 6552 16609 6586 16643
rect 6586 16609 6604 16643
rect 6552 16600 6604 16609
rect 8116 16668 8168 16720
rect 9680 16736 9732 16788
rect 10600 16736 10652 16788
rect 10416 16668 10468 16720
rect 10692 16668 10744 16720
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 5724 16532 5776 16584
rect 8484 16532 8536 16584
rect 8116 16464 8168 16516
rect 9128 16532 9180 16584
rect 9864 16600 9916 16652
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10232 16643 10284 16652
rect 10232 16609 10241 16643
rect 10241 16609 10275 16643
rect 10275 16609 10284 16643
rect 10232 16600 10284 16609
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 12992 16736 13044 16788
rect 12348 16668 12400 16720
rect 12256 16600 12308 16652
rect 5172 16439 5224 16448
rect 5172 16405 5181 16439
rect 5181 16405 5215 16439
rect 5215 16405 5224 16439
rect 5172 16396 5224 16405
rect 7840 16396 7892 16448
rect 8484 16439 8536 16448
rect 8484 16405 8493 16439
rect 8493 16405 8527 16439
rect 8527 16405 8536 16439
rect 8484 16396 8536 16405
rect 9496 16464 9548 16516
rect 9680 16464 9732 16516
rect 11060 16464 11112 16516
rect 9956 16396 10008 16448
rect 10692 16396 10744 16448
rect 10968 16439 11020 16448
rect 10968 16405 10977 16439
rect 10977 16405 11011 16439
rect 11011 16405 11020 16439
rect 10968 16396 11020 16405
rect 12072 16396 12124 16448
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 5172 16192 5224 16244
rect 6000 16192 6052 16244
rect 6552 16192 6604 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 9864 16192 9916 16244
rect 4988 16124 5040 16176
rect 8484 16056 8536 16108
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 10968 16124 11020 16176
rect 11060 16124 11112 16176
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 9036 16056 9088 16108
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 9588 16056 9640 16108
rect 5540 15963 5592 15972
rect 5540 15929 5567 15963
rect 5567 15929 5592 15963
rect 5540 15920 5592 15929
rect 5724 15963 5776 15972
rect 5724 15929 5733 15963
rect 5733 15929 5767 15963
rect 5767 15929 5776 15963
rect 5724 15920 5776 15929
rect 4804 15852 4856 15904
rect 6368 15852 6420 15904
rect 8208 15920 8260 15972
rect 9312 16031 9364 16040
rect 9312 15997 9320 16031
rect 9320 15997 9354 16031
rect 9354 15997 9364 16031
rect 9312 15988 9364 15997
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10968 15988 11020 16040
rect 8668 15852 8720 15904
rect 9128 15852 9180 15904
rect 9404 15852 9456 15904
rect 9680 15852 9732 15904
rect 10416 15852 10468 15904
rect 11612 16031 11664 16040
rect 11612 15997 11621 16031
rect 11621 15997 11655 16031
rect 11655 15997 11664 16031
rect 11612 15988 11664 15997
rect 16120 16192 16172 16244
rect 11796 15988 11848 16040
rect 11520 15963 11572 15972
rect 11520 15929 11529 15963
rect 11529 15929 11563 15963
rect 11563 15929 11572 15963
rect 11520 15920 11572 15929
rect 12072 15988 12124 16040
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 12532 15920 12584 15972
rect 13084 15852 13136 15904
rect 13544 15895 13596 15904
rect 13544 15861 13553 15895
rect 13553 15861 13587 15895
rect 13587 15861 13596 15895
rect 13544 15852 13596 15861
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 5908 15648 5960 15700
rect 4988 15580 5040 15632
rect 6000 15623 6052 15632
rect 6000 15589 6009 15623
rect 6009 15589 6043 15623
rect 6043 15589 6052 15623
rect 6000 15580 6052 15589
rect 8484 15648 8536 15700
rect 10232 15648 10284 15700
rect 2320 15555 2372 15564
rect 2320 15521 2329 15555
rect 2329 15521 2363 15555
rect 2363 15521 2372 15555
rect 2320 15512 2372 15521
rect 3332 15512 3384 15564
rect 4344 15512 4396 15564
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 8116 15512 8168 15564
rect 9036 15555 9088 15564
rect 9036 15521 9045 15555
rect 9045 15521 9079 15555
rect 9079 15521 9088 15555
rect 9036 15512 9088 15521
rect 9128 15555 9180 15564
rect 9128 15521 9138 15555
rect 9138 15521 9172 15555
rect 9172 15521 9180 15555
rect 9128 15512 9180 15521
rect 9312 15555 9364 15564
rect 9312 15521 9321 15555
rect 9321 15521 9355 15555
rect 9355 15521 9364 15555
rect 9312 15512 9364 15521
rect 3424 15376 3476 15428
rect 8576 15487 8628 15496
rect 8576 15453 8585 15487
rect 8585 15453 8619 15487
rect 8619 15453 8628 15487
rect 8576 15444 8628 15453
rect 8668 15444 8720 15496
rect 9220 15444 9272 15496
rect 9588 15512 9640 15564
rect 10416 15580 10468 15632
rect 10968 15691 11020 15700
rect 10968 15657 10977 15691
rect 10977 15657 11011 15691
rect 11011 15657 11020 15691
rect 10968 15648 11020 15657
rect 11520 15648 11572 15700
rect 10232 15555 10284 15564
rect 10232 15521 10241 15555
rect 10241 15521 10275 15555
rect 10275 15521 10284 15555
rect 10232 15512 10284 15521
rect 10508 15512 10560 15564
rect 11244 15512 11296 15564
rect 13084 15555 13136 15564
rect 13084 15521 13093 15555
rect 13093 15521 13127 15555
rect 13127 15521 13136 15555
rect 13084 15512 13136 15521
rect 8024 15376 8076 15428
rect 11336 15376 11388 15428
rect 4344 15308 4396 15360
rect 6000 15308 6052 15360
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7380 15308 7432 15317
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 12072 15308 12124 15360
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 3332 15104 3384 15156
rect 6092 15104 6144 15156
rect 6644 15104 6696 15156
rect 6276 14968 6328 15020
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 3424 14943 3476 14952
rect 3424 14909 3433 14943
rect 3433 14909 3467 14943
rect 3467 14909 3476 14943
rect 3424 14900 3476 14909
rect 4620 14900 4672 14952
rect 4712 14943 4764 14952
rect 4712 14909 4721 14943
rect 4721 14909 4755 14943
rect 4755 14909 4764 14943
rect 4712 14900 4764 14909
rect 7380 14900 7432 14952
rect 8576 14943 8628 14952
rect 7380 14764 7432 14816
rect 8576 14909 8585 14943
rect 8585 14909 8619 14943
rect 8619 14909 8628 14943
rect 8576 14900 8628 14909
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 11796 14943 11848 14952
rect 11796 14909 11805 14943
rect 11805 14909 11839 14943
rect 11839 14909 11848 14943
rect 11796 14900 11848 14909
rect 12532 14968 12584 15020
rect 13084 14900 13136 14952
rect 13820 14900 13872 14952
rect 11152 14832 11204 14884
rect 8208 14764 8260 14816
rect 9772 14764 9824 14816
rect 10232 14764 10284 14816
rect 11704 14764 11756 14816
rect 13912 14764 13964 14816
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 2320 14492 2372 14544
rect 3424 14492 3476 14544
rect 3608 14560 3660 14612
rect 4252 14560 4304 14612
rect 4712 14560 4764 14612
rect 4620 14492 4672 14544
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 13636 14560 13688 14612
rect 8208 14492 8260 14544
rect 2136 14467 2188 14476
rect 2136 14433 2170 14467
rect 2170 14433 2188 14467
rect 2136 14424 2188 14433
rect 3240 14424 3292 14476
rect 5908 14424 5960 14476
rect 6368 14467 6420 14476
rect 6368 14433 6377 14467
rect 6377 14433 6411 14467
rect 6411 14433 6420 14467
rect 6368 14424 6420 14433
rect 6460 14424 6512 14476
rect 4436 14356 4488 14408
rect 7288 14356 7340 14408
rect 7932 14424 7984 14476
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 8024 14356 8076 14408
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 8944 14288 8996 14340
rect 9404 14399 9456 14408
rect 9404 14365 9413 14399
rect 9413 14365 9447 14399
rect 9447 14365 9456 14399
rect 9404 14356 9456 14365
rect 10324 14424 10376 14476
rect 13084 14492 13136 14544
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 11336 14424 11388 14476
rect 12532 14424 12584 14476
rect 13360 14467 13412 14476
rect 13360 14433 13369 14467
rect 13369 14433 13403 14467
rect 13403 14433 13412 14467
rect 13360 14424 13412 14433
rect 13912 14467 13964 14476
rect 13912 14433 13946 14467
rect 13946 14433 13964 14467
rect 13912 14424 13964 14433
rect 12072 14356 12124 14408
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 9220 14220 9272 14272
rect 10784 14220 10836 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 14924 14288 14976 14340
rect 13912 14220 13964 14272
rect 14004 14220 14056 14272
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 2136 14016 2188 14068
rect 3608 13948 3660 14000
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 7288 14059 7340 14068
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7932 14059 7984 14068
rect 7932 14025 7941 14059
rect 7941 14025 7975 14059
rect 7975 14025 7984 14059
rect 7932 14016 7984 14025
rect 8024 14016 8076 14068
rect 5448 13948 5500 14000
rect 3792 13880 3844 13932
rect 4344 13880 4396 13932
rect 9404 14016 9456 14068
rect 13820 14016 13872 14068
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 8668 13948 8720 14000
rect 11336 13991 11388 14000
rect 11336 13957 11345 13991
rect 11345 13957 11379 13991
rect 11379 13957 11388 13991
rect 11336 13948 11388 13957
rect 11428 13948 11480 14000
rect 3240 13855 3292 13864
rect 3240 13821 3249 13855
rect 3249 13821 3283 13855
rect 3283 13821 3292 13855
rect 3240 13812 3292 13821
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 4160 13812 4212 13864
rect 6184 13812 6236 13864
rect 6644 13812 6696 13864
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 5540 13744 5592 13796
rect 5908 13787 5960 13796
rect 5908 13753 5917 13787
rect 5917 13753 5951 13787
rect 5951 13753 5960 13787
rect 5908 13744 5960 13753
rect 7104 13744 7156 13796
rect 8300 13812 8352 13864
rect 8484 13812 8536 13864
rect 12072 13880 12124 13932
rect 13636 13948 13688 14000
rect 12900 13880 12952 13932
rect 13452 13880 13504 13932
rect 8944 13787 8996 13796
rect 4988 13719 5040 13728
rect 4988 13685 4997 13719
rect 4997 13685 5031 13719
rect 5031 13685 5040 13719
rect 4988 13676 5040 13685
rect 6552 13676 6604 13728
rect 6920 13676 6972 13728
rect 8944 13753 8978 13787
rect 8978 13753 8996 13787
rect 8944 13744 8996 13753
rect 11244 13744 11296 13796
rect 11520 13787 11572 13796
rect 11520 13753 11529 13787
rect 11529 13753 11563 13787
rect 11563 13753 11572 13787
rect 11520 13744 11572 13753
rect 12808 13812 12860 13864
rect 13360 13812 13412 13864
rect 14004 13880 14056 13932
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 12532 13719 12584 13728
rect 12532 13685 12541 13719
rect 12541 13685 12575 13719
rect 12575 13685 12584 13719
rect 12532 13676 12584 13685
rect 12808 13676 12860 13728
rect 12992 13719 13044 13728
rect 12992 13685 13001 13719
rect 13001 13685 13035 13719
rect 13035 13685 13044 13719
rect 12992 13676 13044 13685
rect 13636 13676 13688 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 3240 13472 3292 13524
rect 4988 13336 5040 13388
rect 5540 13472 5592 13524
rect 6920 13472 6972 13524
rect 12072 13472 12124 13524
rect 12808 13472 12860 13524
rect 14464 13472 14516 13524
rect 6460 13404 6512 13456
rect 6644 13404 6696 13456
rect 6736 13404 6788 13456
rect 9864 13404 9916 13456
rect 2504 13132 2556 13184
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 5448 13336 5500 13388
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 4804 13175 4856 13184
rect 4804 13141 4813 13175
rect 4813 13141 4847 13175
rect 4847 13141 4856 13175
rect 4804 13132 4856 13141
rect 5908 13268 5960 13320
rect 7104 13336 7156 13388
rect 5908 13132 5960 13184
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 7104 13200 7156 13252
rect 8208 13336 8260 13388
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 9956 13336 10008 13388
rect 12624 13336 12676 13388
rect 13176 13336 13228 13388
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 13728 13379 13780 13388
rect 13728 13345 13737 13379
rect 13737 13345 13771 13379
rect 13771 13345 13780 13379
rect 13728 13336 13780 13345
rect 13912 13336 13964 13388
rect 9772 13268 9824 13320
rect 10048 13268 10100 13320
rect 10600 13268 10652 13320
rect 10232 13132 10284 13184
rect 10968 13132 11020 13184
rect 16672 13132 16724 13184
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 5448 12928 5500 12980
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 9404 12928 9456 12980
rect 9772 12860 9824 12912
rect 2320 12792 2372 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 6736 12792 6788 12844
rect 10140 12928 10192 12980
rect 10324 12903 10376 12912
rect 10324 12869 10333 12903
rect 10333 12869 10367 12903
rect 10367 12869 10376 12903
rect 10324 12860 10376 12869
rect 4620 12724 4672 12776
rect 6184 12724 6236 12776
rect 4252 12656 4304 12708
rect 6920 12724 6972 12776
rect 9956 12724 10008 12776
rect 10048 12767 10100 12776
rect 10048 12733 10060 12767
rect 10060 12733 10094 12767
rect 10094 12733 10100 12767
rect 10048 12724 10100 12733
rect 10232 12724 10284 12776
rect 11520 12928 11572 12980
rect 11612 12928 11664 12980
rect 10692 12903 10744 12912
rect 10692 12869 10701 12903
rect 10701 12869 10735 12903
rect 10735 12869 10744 12903
rect 10692 12860 10744 12869
rect 11796 12903 11848 12912
rect 11796 12869 11805 12903
rect 11805 12869 11839 12903
rect 11839 12869 11848 12903
rect 11796 12860 11848 12869
rect 11980 12860 12032 12912
rect 12348 12860 12400 12912
rect 15108 12860 15160 12912
rect 12532 12792 12584 12844
rect 7288 12656 7340 12708
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 5816 12588 5868 12597
rect 6184 12588 6236 12640
rect 6644 12588 6696 12640
rect 9496 12656 9548 12708
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 12440 12767 12492 12776
rect 12440 12733 12449 12767
rect 12449 12733 12483 12767
rect 12483 12733 12492 12767
rect 12440 12724 12492 12733
rect 13084 12767 13136 12776
rect 13084 12733 13093 12767
rect 13093 12733 13127 12767
rect 13127 12733 13136 12767
rect 13084 12724 13136 12733
rect 13820 12724 13872 12776
rect 10968 12656 11020 12708
rect 13544 12656 13596 12708
rect 10416 12588 10468 12640
rect 10600 12588 10652 12640
rect 10784 12588 10836 12640
rect 11704 12588 11756 12640
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 4160 12384 4212 12436
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 6920 12384 6972 12436
rect 7288 12427 7340 12436
rect 7288 12393 7297 12427
rect 7297 12393 7331 12427
rect 7331 12393 7340 12427
rect 7288 12384 7340 12393
rect 11152 12427 11204 12436
rect 11152 12393 11161 12427
rect 11161 12393 11195 12427
rect 11195 12393 11204 12427
rect 11152 12384 11204 12393
rect 10784 12316 10836 12368
rect 10968 12359 11020 12368
rect 10968 12325 10977 12359
rect 10977 12325 11011 12359
rect 11011 12325 11020 12359
rect 10968 12316 11020 12325
rect 2320 12248 2372 12300
rect 2504 12291 2556 12300
rect 2504 12257 2538 12291
rect 2538 12257 2556 12291
rect 2504 12248 2556 12257
rect 4804 12248 4856 12300
rect 5724 12248 5776 12300
rect 7104 12248 7156 12300
rect 10600 12291 10652 12300
rect 10600 12257 10609 12291
rect 10609 12257 10643 12291
rect 10643 12257 10652 12291
rect 10600 12248 10652 12257
rect 11520 12384 11572 12436
rect 12440 12384 12492 12436
rect 13820 12427 13872 12436
rect 13820 12393 13829 12427
rect 13829 12393 13863 12427
rect 13863 12393 13872 12427
rect 13820 12384 13872 12393
rect 12624 12359 12676 12368
rect 12624 12325 12633 12359
rect 12633 12325 12667 12359
rect 12667 12325 12676 12359
rect 12624 12316 12676 12325
rect 14464 12384 14516 12436
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 12992 12248 13044 12300
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 12716 12223 12768 12232
rect 12716 12189 12725 12223
rect 12725 12189 12759 12223
rect 12759 12189 12768 12223
rect 12716 12180 12768 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 6828 12112 6880 12164
rect 13820 12112 13872 12164
rect 14004 12112 14056 12164
rect 6736 12044 6788 12096
rect 10232 12044 10284 12096
rect 10968 12087 11020 12096
rect 10968 12053 10977 12087
rect 10977 12053 11011 12087
rect 11011 12053 11020 12087
rect 10968 12044 11020 12053
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 5724 11883 5776 11892
rect 5724 11849 5733 11883
rect 5733 11849 5767 11883
rect 5767 11849 5776 11883
rect 5724 11840 5776 11849
rect 6092 11883 6144 11892
rect 6092 11849 6101 11883
rect 6101 11849 6135 11883
rect 6135 11849 6144 11883
rect 6092 11840 6144 11849
rect 10600 11840 10652 11892
rect 13268 11840 13320 11892
rect 13452 11840 13504 11892
rect 10324 11772 10376 11824
rect 10692 11772 10744 11824
rect 12072 11772 12124 11824
rect 6736 11704 6788 11756
rect 12440 11704 12492 11756
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 6184 11679 6236 11688
rect 6184 11645 6193 11679
rect 6193 11645 6227 11679
rect 6227 11645 6236 11679
rect 6184 11636 6236 11645
rect 5448 11568 5500 11620
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 10324 11636 10376 11688
rect 12624 11636 12676 11688
rect 6920 11568 6972 11620
rect 11796 11568 11848 11620
rect 12256 11568 12308 11620
rect 13176 11636 13228 11688
rect 13268 11636 13320 11688
rect 12532 11500 12584 11552
rect 13452 11568 13504 11620
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 14280 11636 14332 11688
rect 14464 11568 14516 11620
rect 14372 11500 14424 11552
rect 14924 11500 14976 11552
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 6828 11296 6880 11348
rect 10048 11339 10100 11348
rect 10048 11305 10057 11339
rect 10057 11305 10091 11339
rect 10091 11305 10100 11339
rect 10048 11296 10100 11305
rect 10324 11296 10376 11348
rect 10876 11296 10928 11348
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 3792 11160 3844 11212
rect 3976 11160 4028 11212
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 8760 11203 8812 11212
rect 8760 11169 8794 11203
rect 8794 11169 8812 11203
rect 8760 11160 8812 11169
rect 11244 11228 11296 11280
rect 11796 11228 11848 11280
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 11060 11160 11112 11212
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 13728 11296 13780 11348
rect 14004 11339 14056 11348
rect 14004 11305 14013 11339
rect 14013 11305 14047 11339
rect 14047 11305 14056 11339
rect 14004 11296 14056 11305
rect 14464 11296 14516 11348
rect 15844 11228 15896 11280
rect 13820 11203 13872 11212
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 14372 11203 14424 11212
rect 14372 11169 14381 11203
rect 14381 11169 14415 11203
rect 14415 11169 14424 11203
rect 14372 11160 14424 11169
rect 14280 11092 14332 11144
rect 9496 11024 9548 11076
rect 9864 10999 9916 11008
rect 9864 10965 9873 10999
rect 9873 10965 9907 10999
rect 9907 10965 9916 10999
rect 9864 10956 9916 10965
rect 10324 10956 10376 11008
rect 10876 10956 10928 11008
rect 11428 10956 11480 11008
rect 12256 10956 12308 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 3976 10752 4028 10804
rect 4988 10752 5040 10804
rect 3792 10684 3844 10736
rect 6184 10684 6236 10736
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 8760 10752 8812 10804
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 8484 10684 8536 10736
rect 4528 10659 4580 10668
rect 4528 10625 4537 10659
rect 4537 10625 4571 10659
rect 4571 10625 4580 10659
rect 4528 10616 4580 10625
rect 4988 10659 5040 10668
rect 4988 10625 4997 10659
rect 4997 10625 5031 10659
rect 5031 10625 5040 10659
rect 4988 10616 5040 10625
rect 7656 10616 7708 10668
rect 10048 10616 10100 10668
rect 3976 10548 4028 10600
rect 4620 10591 4672 10600
rect 4620 10557 4629 10591
rect 4629 10557 4663 10591
rect 4663 10557 4672 10591
rect 4620 10548 4672 10557
rect 5540 10548 5592 10600
rect 6644 10548 6696 10600
rect 6736 10591 6788 10600
rect 6736 10557 6748 10591
rect 6748 10557 6782 10591
rect 6782 10557 6788 10591
rect 6736 10548 6788 10557
rect 7104 10548 7156 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 7472 10591 7524 10600
rect 7472 10557 7481 10591
rect 7481 10557 7515 10591
rect 7515 10557 7524 10591
rect 7472 10548 7524 10557
rect 9404 10548 9456 10600
rect 10416 10591 10468 10600
rect 10416 10557 10425 10591
rect 10425 10557 10459 10591
rect 10459 10557 10468 10591
rect 10416 10548 10468 10557
rect 6368 10480 6420 10532
rect 4804 10412 4856 10464
rect 5448 10412 5500 10464
rect 10508 10480 10560 10532
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 10876 10548 10928 10557
rect 13176 10616 13228 10668
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15292 10616 15344 10625
rect 16212 10616 16264 10668
rect 7012 10412 7064 10464
rect 8024 10412 8076 10464
rect 9864 10412 9916 10464
rect 10968 10412 11020 10464
rect 15016 10548 15068 10600
rect 15384 10548 15436 10600
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 11888 10412 11940 10464
rect 12992 10412 13044 10464
rect 13728 10412 13780 10464
rect 16028 10412 16080 10464
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 3792 10251 3844 10260
rect 3792 10217 3817 10251
rect 3817 10217 3844 10251
rect 3792 10208 3844 10217
rect 3976 10251 4028 10260
rect 3976 10217 3985 10251
rect 3985 10217 4019 10251
rect 4019 10217 4028 10251
rect 3976 10208 4028 10217
rect 4252 10115 4304 10124
rect 4252 10081 4264 10115
rect 4264 10081 4298 10115
rect 4298 10081 4304 10115
rect 4252 10072 4304 10081
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 4436 10072 4488 10124
rect 6736 10251 6788 10260
rect 6736 10217 6745 10251
rect 6745 10217 6779 10251
rect 6779 10217 6788 10251
rect 6736 10208 6788 10217
rect 5356 10115 5408 10124
rect 5356 10081 5365 10115
rect 5365 10081 5399 10115
rect 5399 10081 5408 10115
rect 5356 10072 5408 10081
rect 7380 10208 7432 10260
rect 7472 10251 7524 10260
rect 7472 10217 7481 10251
rect 7481 10217 7515 10251
rect 7515 10217 7524 10251
rect 7472 10208 7524 10217
rect 7656 10251 7708 10260
rect 7656 10217 7665 10251
rect 7665 10217 7699 10251
rect 7699 10217 7708 10251
rect 7656 10208 7708 10217
rect 8300 10208 8352 10260
rect 12072 10208 12124 10260
rect 13452 10208 13504 10260
rect 6184 10004 6236 10056
rect 4436 9936 4488 9988
rect 5080 9936 5132 9988
rect 5448 9979 5500 9988
rect 5448 9945 5457 9979
rect 5457 9945 5491 9979
rect 5491 9945 5500 9979
rect 5448 9936 5500 9945
rect 5540 9936 5592 9988
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 8392 10140 8444 10192
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 8208 10115 8260 10124
rect 8208 10081 8217 10115
rect 8217 10081 8251 10115
rect 8251 10081 8260 10115
rect 8208 10072 8260 10081
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 3884 9868 3936 9920
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 6828 9868 6880 9920
rect 8760 10004 8812 10056
rect 9404 10072 9456 10124
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11428 10115 11480 10124
rect 11428 10081 11437 10115
rect 11437 10081 11471 10115
rect 11471 10081 11480 10115
rect 11428 10072 11480 10081
rect 11520 10072 11572 10124
rect 12716 10140 12768 10192
rect 12072 10004 12124 10056
rect 8024 9936 8076 9988
rect 13084 10115 13136 10124
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 13268 10047 13320 10056
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 14096 10072 14148 10124
rect 14832 10115 14884 10124
rect 14832 10081 14836 10115
rect 14836 10081 14870 10115
rect 14870 10081 14884 10115
rect 14832 10072 14884 10081
rect 13912 10004 13964 10056
rect 14372 10004 14424 10056
rect 13176 9868 13228 9920
rect 13728 9868 13780 9920
rect 13820 9911 13872 9920
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 14004 9868 14056 9920
rect 15200 10115 15252 10124
rect 15200 10081 15208 10115
rect 15208 10081 15242 10115
rect 15242 10081 15252 10115
rect 15200 10072 15252 10081
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 15476 10140 15528 10192
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 16488 10072 16540 10124
rect 15568 9868 15620 9920
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 4528 9664 4580 9716
rect 5632 9664 5684 9716
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 6460 9664 6512 9716
rect 7196 9707 7248 9716
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 12072 9664 12124 9716
rect 12440 9664 12492 9716
rect 13176 9664 13228 9716
rect 13268 9664 13320 9716
rect 14832 9664 14884 9716
rect 5448 9596 5500 9648
rect 4712 9528 4764 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 6920 9596 6972 9648
rect 8208 9596 8260 9648
rect 9680 9596 9732 9648
rect 11612 9596 11664 9648
rect 5080 9528 5132 9537
rect 4344 9392 4396 9444
rect 5816 9460 5868 9512
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6736 9528 6788 9580
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 7012 9528 7064 9580
rect 8024 9528 8076 9580
rect 7656 9503 7708 9512
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 9404 9528 9456 9580
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 11060 9503 11112 9512
rect 11060 9469 11069 9503
rect 11069 9469 11103 9503
rect 11103 9469 11112 9503
rect 11060 9460 11112 9469
rect 9496 9392 9548 9444
rect 10876 9392 10928 9444
rect 11612 9503 11664 9512
rect 11612 9469 11621 9503
rect 11621 9469 11655 9503
rect 11655 9469 11664 9503
rect 11612 9460 11664 9469
rect 12256 9528 12308 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12992 9528 13044 9580
rect 13452 9596 13504 9648
rect 15200 9596 15252 9648
rect 15660 9596 15712 9648
rect 15844 9639 15896 9648
rect 15844 9605 15853 9639
rect 15853 9605 15887 9639
rect 15887 9605 15896 9639
rect 15844 9596 15896 9605
rect 12348 9503 12400 9512
rect 12348 9469 12353 9503
rect 12353 9469 12387 9503
rect 12387 9469 12400 9503
rect 12348 9460 12400 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 12072 9392 12124 9444
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 14004 9503 14056 9512
rect 14004 9469 14039 9503
rect 14039 9469 14056 9503
rect 14004 9460 14056 9469
rect 14188 9503 14240 9512
rect 14188 9469 14197 9503
rect 14197 9469 14231 9503
rect 14231 9469 14240 9503
rect 14188 9460 14240 9469
rect 14464 9460 14516 9512
rect 14372 9392 14424 9444
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 16028 9528 16080 9580
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16212 9503 16264 9512
rect 16212 9469 16221 9503
rect 16221 9469 16255 9503
rect 16255 9469 16264 9503
rect 16212 9460 16264 9469
rect 6000 9324 6052 9376
rect 6276 9324 6328 9376
rect 6552 9324 6604 9376
rect 7012 9324 7064 9376
rect 7748 9324 7800 9376
rect 8576 9324 8628 9376
rect 9036 9324 9088 9376
rect 10508 9324 10560 9376
rect 10968 9324 11020 9376
rect 12440 9324 12492 9376
rect 12716 9324 12768 9376
rect 13084 9324 13136 9376
rect 13636 9324 13688 9376
rect 13820 9324 13872 9376
rect 14004 9324 14056 9376
rect 15384 9324 15436 9376
rect 15568 9435 15620 9444
rect 15568 9401 15577 9435
rect 15577 9401 15611 9435
rect 15611 9401 15620 9435
rect 16396 9503 16448 9512
rect 16396 9469 16405 9503
rect 16405 9469 16439 9503
rect 16439 9469 16448 9503
rect 16396 9460 16448 9469
rect 16488 9503 16540 9512
rect 16488 9469 16497 9503
rect 16497 9469 16531 9503
rect 16531 9469 16540 9503
rect 16488 9460 16540 9469
rect 15568 9392 15620 9401
rect 16580 9435 16632 9444
rect 16580 9401 16589 9435
rect 16589 9401 16623 9435
rect 16623 9401 16632 9435
rect 16580 9392 16632 9401
rect 15936 9324 15988 9376
rect 16396 9324 16448 9376
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 6828 9052 6880 9104
rect 7104 9163 7156 9172
rect 7104 9129 7113 9163
rect 7113 9129 7147 9163
rect 7147 9129 7156 9163
rect 7104 9120 7156 9129
rect 7656 9120 7708 9172
rect 8116 9120 8168 9172
rect 6552 8984 6604 9036
rect 7288 9052 7340 9104
rect 7748 9052 7800 9104
rect 7564 9027 7616 9036
rect 7564 8993 7573 9027
rect 7573 8993 7607 9027
rect 7607 8993 7616 9027
rect 7564 8984 7616 8993
rect 7840 9027 7892 9036
rect 7840 8993 7849 9027
rect 7849 8993 7883 9027
rect 7883 8993 7892 9027
rect 7840 8984 7892 8993
rect 7932 8848 7984 8900
rect 8576 9095 8628 9104
rect 8576 9061 8585 9095
rect 8585 9061 8619 9095
rect 8619 9061 8628 9095
rect 8576 9052 8628 9061
rect 8668 9052 8720 9104
rect 9128 9052 9180 9104
rect 10140 9120 10192 9172
rect 10324 9120 10376 9172
rect 11428 9120 11480 9172
rect 8760 9027 8812 9036
rect 8760 8993 8769 9027
rect 8769 8993 8803 9027
rect 8803 8993 8812 9027
rect 8760 8984 8812 8993
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 9588 9027 9640 9036
rect 9588 8993 9597 9027
rect 9597 8993 9631 9027
rect 9631 8993 9640 9027
rect 9588 8984 9640 8993
rect 8668 8916 8720 8968
rect 8944 8916 8996 8968
rect 9220 8916 9272 8968
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 10968 8984 11020 9036
rect 11520 9027 11572 9036
rect 11520 8993 11529 9027
rect 11529 8993 11563 9027
rect 11563 8993 11572 9027
rect 11520 8984 11572 8993
rect 11980 8984 12032 9036
rect 12716 9120 12768 9172
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 10232 8916 10284 8968
rect 12440 8916 12492 8968
rect 9956 8848 10008 8900
rect 10416 8848 10468 8900
rect 11060 8848 11112 8900
rect 5448 8780 5500 8832
rect 5908 8780 5960 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7380 8780 7432 8832
rect 8024 8780 8076 8832
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 9036 8823 9088 8832
rect 9036 8789 9057 8823
rect 9057 8789 9088 8823
rect 9036 8780 9088 8789
rect 9772 8780 9824 8832
rect 11244 8780 11296 8832
rect 12624 8780 12676 8832
rect 12992 8916 13044 8968
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 14188 9120 14240 9172
rect 14372 9120 14424 9172
rect 16580 9120 16632 9172
rect 13360 8916 13412 8968
rect 13728 8984 13780 9036
rect 14096 9027 14148 9036
rect 14096 8993 14105 9027
rect 14105 8993 14139 9027
rect 14139 8993 14148 9027
rect 14096 8984 14148 8993
rect 14924 8984 14976 9036
rect 15384 9027 15436 9036
rect 15384 8993 15393 9027
rect 15393 8993 15427 9027
rect 15427 8993 15436 9027
rect 15384 8984 15436 8993
rect 13636 8916 13688 8968
rect 15016 8916 15068 8968
rect 16212 8984 16264 9036
rect 15936 8916 15988 8968
rect 16580 8984 16632 9036
rect 17224 8984 17276 9036
rect 14464 8848 14516 8900
rect 16580 8848 16632 8900
rect 13084 8780 13136 8832
rect 13820 8780 13872 8832
rect 14280 8823 14332 8832
rect 14280 8789 14289 8823
rect 14289 8789 14323 8823
rect 14323 8789 14332 8823
rect 14280 8780 14332 8789
rect 15568 8780 15620 8832
rect 16120 8780 16172 8832
rect 16396 8780 16448 8832
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 4620 8576 4672 8628
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 9496 8576 9548 8628
rect 10140 8576 10192 8628
rect 10600 8576 10652 8628
rect 11428 8576 11480 8628
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 4068 8508 4120 8560
rect 3792 8415 3844 8424
rect 3792 8381 3801 8415
rect 3801 8381 3835 8415
rect 3835 8381 3844 8415
rect 3792 8372 3844 8381
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 4528 8440 4580 8492
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 4988 8440 5040 8492
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 4712 8236 4764 8288
rect 5632 8304 5684 8356
rect 6092 8372 6144 8424
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 6736 8440 6788 8492
rect 7840 8440 7892 8492
rect 6460 8372 6512 8424
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 7012 8372 7064 8424
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 7932 8372 7984 8424
rect 9772 8508 9824 8560
rect 9956 8508 10008 8560
rect 10140 8440 10192 8492
rect 10508 8508 10560 8560
rect 10876 8551 10928 8560
rect 10876 8517 10885 8551
rect 10885 8517 10919 8551
rect 10919 8517 10928 8551
rect 10876 8508 10928 8517
rect 10968 8551 11020 8560
rect 10968 8517 10977 8551
rect 10977 8517 11011 8551
rect 11011 8517 11020 8551
rect 10968 8508 11020 8517
rect 12624 8508 12676 8560
rect 13452 8508 13504 8560
rect 14924 8576 14976 8628
rect 15568 8576 15620 8628
rect 16212 8576 16264 8628
rect 17224 8576 17276 8628
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 9956 8372 10008 8424
rect 10416 8372 10468 8424
rect 10600 8372 10652 8424
rect 8944 8347 8996 8356
rect 8944 8313 8953 8347
rect 8953 8313 8987 8347
rect 8987 8313 8996 8347
rect 8944 8304 8996 8313
rect 9496 8304 9548 8356
rect 6276 8236 6328 8288
rect 7104 8279 7156 8288
rect 7104 8245 7113 8279
rect 7113 8245 7147 8279
rect 7147 8245 7156 8279
rect 7104 8236 7156 8245
rect 8300 8236 8352 8288
rect 10232 8304 10284 8356
rect 10048 8236 10100 8288
rect 11060 8304 11112 8356
rect 11428 8304 11480 8356
rect 13268 8440 13320 8492
rect 11888 8372 11940 8424
rect 14280 8508 14332 8560
rect 14188 8415 14240 8424
rect 14188 8381 14197 8415
rect 14197 8381 14231 8415
rect 14231 8381 14240 8415
rect 14188 8372 14240 8381
rect 14280 8372 14332 8424
rect 16028 8440 16080 8492
rect 10784 8236 10836 8288
rect 11612 8236 11664 8288
rect 13912 8347 13964 8356
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 14004 8347 14056 8356
rect 14004 8313 14039 8347
rect 14039 8313 14056 8347
rect 14004 8304 14056 8313
rect 14464 8304 14516 8356
rect 15384 8372 15436 8424
rect 16764 8372 16816 8424
rect 16396 8347 16448 8356
rect 16396 8313 16405 8347
rect 16405 8313 16439 8347
rect 16439 8313 16448 8347
rect 16396 8304 16448 8313
rect 15476 8236 15528 8288
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 4252 8032 4304 8084
rect 4988 8032 5040 8084
rect 6368 8032 6420 8084
rect 7196 8032 7248 8084
rect 9588 8032 9640 8084
rect 10140 8075 10192 8084
rect 10140 8041 10167 8075
rect 10167 8041 10192 8075
rect 10140 8032 10192 8041
rect 10968 8032 11020 8084
rect 11980 8032 12032 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 13912 8032 13964 8084
rect 16212 8032 16264 8084
rect 16764 8032 16816 8084
rect 3424 7939 3476 7948
rect 3424 7905 3442 7939
rect 3442 7905 3476 7939
rect 3424 7896 3476 7905
rect 3976 7896 4028 7948
rect 3792 7828 3844 7880
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 4804 7828 4856 7880
rect 4988 7939 5040 7948
rect 4988 7905 4997 7939
rect 4997 7905 5031 7939
rect 5031 7905 5040 7939
rect 4988 7896 5040 7905
rect 5632 7896 5684 7948
rect 5724 7896 5776 7948
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 9496 7964 9548 8016
rect 10876 7964 10928 8016
rect 12808 7964 12860 8016
rect 6736 7896 6788 7948
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 10140 7896 10192 7948
rect 16580 7964 16632 8016
rect 17224 8007 17276 8016
rect 17224 7973 17233 8007
rect 17233 7973 17267 8007
rect 17267 7973 17276 8007
rect 17224 7964 17276 7973
rect 4068 7735 4120 7744
rect 4068 7701 4077 7735
rect 4077 7701 4111 7735
rect 4111 7701 4120 7735
rect 4068 7692 4120 7701
rect 4344 7735 4396 7744
rect 4344 7701 4353 7735
rect 4353 7701 4387 7735
rect 4387 7701 4396 7735
rect 4344 7692 4396 7701
rect 6644 7692 6696 7744
rect 7932 7692 7984 7744
rect 10232 7760 10284 7812
rect 10508 7692 10560 7744
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 12624 7760 12676 7812
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 13820 7896 13872 7948
rect 15016 7896 15068 7948
rect 15200 7939 15252 7948
rect 15200 7905 15209 7939
rect 15209 7905 15243 7939
rect 15243 7905 15252 7939
rect 15200 7896 15252 7905
rect 15384 7939 15436 7948
rect 15384 7905 15393 7939
rect 15393 7905 15427 7939
rect 15427 7905 15436 7939
rect 15384 7896 15436 7905
rect 13544 7828 13596 7880
rect 15568 7896 15620 7948
rect 15752 7939 15804 7948
rect 15752 7905 15761 7939
rect 15761 7905 15795 7939
rect 15795 7905 15804 7939
rect 15752 7896 15804 7905
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 16304 7939 16356 7948
rect 16304 7905 16308 7939
rect 16308 7905 16342 7939
rect 16342 7905 16356 7939
rect 16304 7896 16356 7905
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 14372 7760 14424 7812
rect 14004 7692 14056 7744
rect 15936 7735 15988 7744
rect 15936 7701 15945 7735
rect 15945 7701 15979 7735
rect 15979 7701 15988 7735
rect 15936 7692 15988 7701
rect 16580 7828 16632 7880
rect 16764 7939 16816 7948
rect 16764 7905 16773 7939
rect 16773 7905 16807 7939
rect 16807 7905 16816 7939
rect 16764 7896 16816 7905
rect 16764 7760 16816 7812
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 3424 7531 3476 7540
rect 3424 7497 3433 7531
rect 3433 7497 3467 7531
rect 3467 7497 3476 7531
rect 3424 7488 3476 7497
rect 4344 7488 4396 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 6184 7488 6236 7540
rect 6460 7488 6512 7540
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 3884 7284 3936 7336
rect 4160 7284 4212 7336
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 5448 7420 5500 7472
rect 5908 7420 5960 7472
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 7472 7420 7524 7472
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 5540 7352 5592 7404
rect 5540 7216 5592 7268
rect 5724 7284 5776 7336
rect 5908 7284 5960 7336
rect 7104 7284 7156 7336
rect 7932 7352 7984 7404
rect 7196 7216 7248 7268
rect 6460 7148 6512 7200
rect 7104 7148 7156 7200
rect 8392 7531 8444 7540
rect 8392 7497 8401 7531
rect 8401 7497 8435 7531
rect 8435 7497 8444 7531
rect 8392 7488 8444 7497
rect 11980 7488 12032 7540
rect 12900 7488 12952 7540
rect 13636 7488 13688 7540
rect 15752 7488 15804 7540
rect 16488 7488 16540 7540
rect 12808 7420 12860 7472
rect 8300 7352 8352 7404
rect 8208 7284 8260 7336
rect 11520 7352 11572 7404
rect 12992 7352 13044 7404
rect 10508 7284 10560 7336
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12256 7327 12308 7336
rect 12256 7293 12265 7327
rect 12265 7293 12299 7327
rect 12299 7293 12308 7327
rect 12256 7284 12308 7293
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 15936 7352 15988 7404
rect 13268 7284 13320 7336
rect 8484 7216 8536 7268
rect 9312 7216 9364 7268
rect 12072 7216 12124 7268
rect 13452 7216 13504 7268
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 15476 7284 15528 7336
rect 16488 7327 16540 7336
rect 16488 7293 16497 7327
rect 16497 7293 16531 7327
rect 16531 7293 16540 7327
rect 16488 7284 16540 7293
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 15200 7259 15252 7268
rect 15200 7225 15209 7259
rect 15209 7225 15243 7259
rect 15243 7225 15252 7259
rect 15200 7216 15252 7225
rect 15384 7216 15436 7268
rect 7656 7148 7708 7200
rect 11980 7148 12032 7200
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 4804 6944 4856 6996
rect 5356 6944 5408 6996
rect 6276 6944 6328 6996
rect 6368 6944 6420 6996
rect 10968 6944 11020 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 12164 6944 12216 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 12900 6944 12952 6996
rect 15476 6944 15528 6996
rect 4804 6808 4856 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 5632 6740 5684 6792
rect 5908 6740 5960 6792
rect 4712 6672 4764 6724
rect 7012 6851 7064 6860
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 8208 6876 8260 6928
rect 10876 6876 10928 6928
rect 7288 6740 7340 6792
rect 8668 6808 8720 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 8208 6740 8260 6792
rect 8576 6783 8628 6792
rect 8576 6749 8585 6783
rect 8585 6749 8619 6783
rect 8619 6749 8628 6783
rect 8576 6740 8628 6749
rect 7932 6672 7984 6724
rect 8024 6672 8076 6724
rect 10416 6672 10468 6724
rect 11428 6672 11480 6724
rect 4068 6604 4120 6656
rect 5080 6604 5132 6656
rect 5540 6604 5592 6656
rect 6000 6604 6052 6656
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 11244 6604 11296 6656
rect 11612 6808 11664 6860
rect 12072 6808 12124 6860
rect 12256 6808 12308 6860
rect 12624 6851 12676 6860
rect 12624 6817 12633 6851
rect 12633 6817 12667 6851
rect 12667 6817 12676 6851
rect 12624 6808 12676 6817
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 13268 6851 13320 6860
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 13820 6808 13872 6860
rect 15660 6808 15712 6860
rect 15936 6808 15988 6860
rect 16396 6808 16448 6860
rect 15384 6783 15436 6792
rect 15384 6749 15393 6783
rect 15393 6749 15427 6783
rect 15427 6749 15436 6783
rect 15384 6740 15436 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 15568 6740 15620 6792
rect 11888 6604 11940 6656
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 14648 6604 14700 6656
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 3608 6400 3660 6452
rect 3792 6264 3844 6316
rect 5448 6400 5500 6452
rect 5264 6332 5316 6384
rect 7104 6400 7156 6452
rect 8208 6400 8260 6452
rect 8944 6400 8996 6452
rect 11612 6443 11664 6452
rect 11612 6409 11621 6443
rect 11621 6409 11655 6443
rect 11655 6409 11664 6443
rect 11612 6400 11664 6409
rect 4804 6196 4856 6248
rect 5080 6239 5132 6248
rect 5080 6205 5089 6239
rect 5089 6205 5123 6239
rect 5123 6205 5132 6239
rect 5080 6196 5132 6205
rect 5724 6264 5776 6316
rect 5356 6196 5408 6248
rect 5448 6196 5500 6248
rect 5908 6307 5960 6316
rect 5908 6273 5917 6307
rect 5917 6273 5951 6307
rect 5951 6273 5960 6307
rect 5908 6264 5960 6273
rect 6736 6264 6788 6316
rect 6000 6239 6052 6248
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 7380 6196 7432 6248
rect 7840 6196 7892 6248
rect 7932 6239 7984 6248
rect 7932 6205 7941 6239
rect 7941 6205 7975 6239
rect 7975 6205 7984 6239
rect 7932 6196 7984 6205
rect 8300 6332 8352 6384
rect 11428 6332 11480 6384
rect 15568 6400 15620 6452
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 12072 6332 12124 6384
rect 8484 6264 8536 6316
rect 9680 6196 9732 6248
rect 13176 6264 13228 6316
rect 14648 6375 14700 6384
rect 14648 6341 14657 6375
rect 14657 6341 14691 6375
rect 14691 6341 14700 6375
rect 14648 6332 14700 6341
rect 6184 6128 6236 6180
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 5540 6060 5592 6069
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 5816 6060 5868 6112
rect 8208 6128 8260 6180
rect 11796 6196 11848 6248
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8024 6060 8076 6112
rect 8484 6060 8536 6112
rect 9404 6060 9456 6112
rect 11244 6128 11296 6180
rect 13544 6239 13596 6248
rect 13544 6205 13553 6239
rect 13553 6205 13587 6239
rect 13587 6205 13596 6239
rect 13544 6196 13596 6205
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 13912 6239 13964 6248
rect 13912 6205 13921 6239
rect 13921 6205 13955 6239
rect 13955 6205 13964 6239
rect 13912 6196 13964 6205
rect 14280 6196 14332 6248
rect 15936 6307 15988 6316
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 16396 6264 16448 6316
rect 15476 6196 15528 6248
rect 11796 6060 11848 6112
rect 13084 6060 13136 6112
rect 13820 6060 13872 6112
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 14280 6060 14332 6112
rect 15016 6128 15068 6180
rect 15292 6128 15344 6180
rect 16028 6239 16080 6248
rect 16028 6205 16037 6239
rect 16037 6205 16071 6239
rect 16071 6205 16080 6239
rect 16028 6196 16080 6205
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 16580 6128 16632 6180
rect 17224 6171 17276 6180
rect 17224 6137 17233 6171
rect 17233 6137 17267 6171
rect 17267 6137 17276 6171
rect 17224 6128 17276 6137
rect 15200 6060 15252 6112
rect 16028 6060 16080 6112
rect 16396 6060 16448 6112
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4068 5720 4120 5772
rect 5632 5856 5684 5908
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 5540 5788 5592 5840
rect 9680 5856 9732 5908
rect 12532 5856 12584 5908
rect 14096 5856 14148 5908
rect 14924 5856 14976 5908
rect 15016 5899 15068 5908
rect 15016 5865 15025 5899
rect 15025 5865 15059 5899
rect 15059 5865 15068 5899
rect 15016 5856 15068 5865
rect 5448 5763 5500 5772
rect 5448 5729 5457 5763
rect 5457 5729 5491 5763
rect 5491 5729 5500 5763
rect 5448 5720 5500 5729
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6000 5763 6052 5772
rect 6000 5729 6007 5763
rect 6007 5729 6052 5763
rect 6000 5720 6052 5729
rect 4988 5652 5040 5704
rect 6184 5652 6236 5704
rect 6828 5763 6880 5772
rect 6828 5729 6837 5763
rect 6837 5729 6871 5763
rect 6871 5729 6880 5763
rect 6828 5720 6880 5729
rect 7196 5720 7248 5772
rect 7380 5763 7432 5772
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 9496 5720 9548 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 13084 5763 13136 5772
rect 13084 5729 13093 5763
rect 13093 5729 13127 5763
rect 13127 5729 13136 5763
rect 13084 5720 13136 5729
rect 13176 5763 13228 5772
rect 13176 5729 13185 5763
rect 13185 5729 13219 5763
rect 13219 5729 13228 5763
rect 13176 5720 13228 5729
rect 14280 5788 14332 5840
rect 13452 5720 13504 5772
rect 14004 5763 14056 5772
rect 14004 5729 14013 5763
rect 14013 5729 14047 5763
rect 14047 5729 14056 5763
rect 14004 5720 14056 5729
rect 7840 5652 7892 5704
rect 8300 5652 8352 5704
rect 8576 5652 8628 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 13268 5652 13320 5704
rect 7380 5584 7432 5636
rect 11888 5584 11940 5636
rect 13820 5584 13872 5636
rect 14464 5720 14516 5772
rect 15016 5720 15068 5772
rect 15660 5720 15712 5772
rect 16028 5720 16080 5772
rect 16396 5763 16448 5772
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 16580 5720 16632 5772
rect 15476 5652 15528 5704
rect 15016 5584 15068 5636
rect 15568 5584 15620 5636
rect 16212 5584 16264 5636
rect 17224 5720 17276 5772
rect 3976 5516 4028 5568
rect 4896 5516 4948 5568
rect 5540 5516 5592 5568
rect 5816 5516 5868 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 7104 5516 7156 5568
rect 9404 5516 9456 5568
rect 11428 5516 11480 5568
rect 14648 5516 14700 5568
rect 14924 5516 14976 5568
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 6460 5312 6512 5364
rect 6644 5312 6696 5364
rect 5080 5244 5132 5296
rect 6552 5176 6604 5228
rect 6920 5108 6972 5160
rect 7288 5108 7340 5160
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11980 5312 12032 5364
rect 12900 5355 12952 5364
rect 12900 5321 12909 5355
rect 12909 5321 12943 5355
rect 12943 5321 12952 5355
rect 12900 5312 12952 5321
rect 13176 5312 13228 5364
rect 15476 5355 15528 5364
rect 15476 5321 15485 5355
rect 15485 5321 15519 5355
rect 15519 5321 15528 5355
rect 15476 5312 15528 5321
rect 16028 5312 16080 5364
rect 7748 5108 7800 5160
rect 8484 5244 8536 5296
rect 8576 5244 8628 5296
rect 11152 5244 11204 5296
rect 12808 5244 12860 5296
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 10876 5176 10928 5228
rect 8484 5108 8536 5160
rect 6000 5040 6052 5092
rect 6644 5040 6696 5092
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 5816 5015 5868 5024
rect 5816 4981 5825 5015
rect 5825 4981 5859 5015
rect 5859 4981 5868 5015
rect 5816 4972 5868 4981
rect 8944 5108 8996 5160
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 12072 5176 12124 5228
rect 12440 5151 12492 5160
rect 12440 5117 12449 5151
rect 12449 5117 12483 5151
rect 12483 5117 12492 5151
rect 12440 5108 12492 5117
rect 14372 5176 14424 5228
rect 7932 4972 7984 5024
rect 8024 4972 8076 5024
rect 11060 5040 11112 5092
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 13820 5108 13872 5160
rect 14188 5151 14240 5160
rect 14188 5117 14197 5151
rect 14197 5117 14231 5151
rect 14231 5117 14240 5151
rect 14188 5108 14240 5117
rect 14924 5219 14976 5228
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 15384 5176 15436 5228
rect 15200 5151 15252 5160
rect 15200 5117 15209 5151
rect 15209 5117 15243 5151
rect 15243 5117 15252 5151
rect 15200 5108 15252 5117
rect 15476 5108 15528 5160
rect 16212 5108 16264 5160
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 16488 5151 16540 5160
rect 16488 5117 16497 5151
rect 16497 5117 16531 5151
rect 16531 5117 16540 5151
rect 16488 5108 16540 5117
rect 11520 4972 11572 5024
rect 12900 4972 12952 5024
rect 13084 5015 13136 5024
rect 13084 4981 13093 5015
rect 13093 4981 13127 5015
rect 13127 4981 13136 5015
rect 13084 4972 13136 4981
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14372 4972 14424 5024
rect 14648 5015 14700 5024
rect 14648 4981 14657 5015
rect 14657 4981 14691 5015
rect 14691 4981 14700 5015
rect 14648 4972 14700 4981
rect 14924 4972 14976 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 6920 4768 6972 4820
rect 6368 4632 6420 4684
rect 7840 4768 7892 4820
rect 7380 4700 7432 4752
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 8576 4700 8628 4752
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 7840 4675 7892 4684
rect 7840 4641 7849 4675
rect 7849 4641 7883 4675
rect 7883 4641 7892 4675
rect 7840 4632 7892 4641
rect 7932 4675 7984 4684
rect 7932 4641 7941 4675
rect 7941 4641 7975 4675
rect 7975 4641 7984 4675
rect 7932 4632 7984 4641
rect 8392 4675 8444 4684
rect 8392 4641 8401 4675
rect 8401 4641 8435 4675
rect 8435 4641 8444 4675
rect 8392 4632 8444 4641
rect 10968 4768 11020 4820
rect 12348 4768 12400 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 12716 4811 12768 4820
rect 12716 4777 12725 4811
rect 12725 4777 12759 4811
rect 12759 4777 12768 4811
rect 12716 4768 12768 4777
rect 12900 4768 12952 4820
rect 14280 4768 14332 4820
rect 14464 4768 14516 4820
rect 10876 4632 10928 4684
rect 11520 4632 11572 4684
rect 11980 4632 12032 4684
rect 13084 4700 13136 4752
rect 12716 4675 12768 4684
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 14096 4632 14148 4684
rect 14280 4632 14332 4684
rect 14556 4675 14608 4684
rect 14556 4641 14565 4675
rect 14565 4641 14599 4675
rect 14599 4641 14608 4675
rect 14556 4632 14608 4641
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 14924 4632 14976 4684
rect 12440 4564 12492 4616
rect 12716 4496 12768 4548
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 8392 4428 8444 4480
rect 8668 4428 8720 4480
rect 12900 4428 12952 4480
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 14004 4607 14056 4616
rect 14004 4573 14013 4607
rect 14013 4573 14047 4607
rect 14047 4573 14056 4607
rect 14004 4564 14056 4573
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 15476 4675 15528 4684
rect 15476 4641 15485 4675
rect 15485 4641 15519 4675
rect 15519 4641 15528 4675
rect 15476 4632 15528 4641
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 16120 4632 16172 4684
rect 13544 4496 13596 4548
rect 13820 4496 13872 4548
rect 14740 4496 14792 4548
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 8668 4267 8720 4276
rect 8668 4233 8677 4267
rect 8677 4233 8711 4267
rect 8711 4233 8720 4267
rect 8668 4224 8720 4233
rect 11980 4224 12032 4276
rect 12900 4224 12952 4276
rect 13728 4224 13780 4276
rect 7380 4156 7432 4208
rect 8944 4156 8996 4208
rect 3976 4020 4028 4072
rect 8300 4020 8352 4072
rect 8392 4063 8444 4072
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 11428 4020 11480 4072
rect 5632 3952 5684 4004
rect 8944 3952 8996 4004
rect 11152 3995 11204 4004
rect 11152 3961 11186 3995
rect 11186 3961 11204 3995
rect 11152 3952 11204 3961
rect 11336 3952 11388 4004
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 13820 4156 13872 4208
rect 14464 4224 14516 4276
rect 14556 4267 14608 4276
rect 14556 4233 14565 4267
rect 14565 4233 14599 4267
rect 14599 4233 14608 4267
rect 14556 4224 14608 4233
rect 16304 4156 16356 4208
rect 13176 4088 13228 4140
rect 13728 4063 13780 4072
rect 13728 4029 13737 4063
rect 13737 4029 13771 4063
rect 13771 4029 13780 4063
rect 13728 4020 13780 4029
rect 14924 4088 14976 4140
rect 15016 4020 15068 4072
rect 14004 3952 14056 4004
rect 7196 3927 7248 3936
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 9680 3884 9732 3936
rect 11520 3884 11572 3936
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 10876 3680 10928 3732
rect 12808 3680 12860 3732
rect 7196 3612 7248 3664
rect 8300 3544 8352 3596
rect 8576 3544 8628 3596
rect 9680 3544 9732 3596
rect 11060 3612 11112 3664
rect 11428 3612 11480 3664
rect 12992 3340 13044 3392
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 3700 2864 3752 2916
rect 6184 2796 6236 2848
rect 11796 2796 11848 2848
rect 12808 2796 12860 2848
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 8668 2592 8720 2644
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 10232 2524 10284 2576
rect 15108 2524 15160 2576
rect 11060 2388 11112 2440
rect 14280 2388 14332 2440
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 11060 1844 11112 1896
rect 10600 1776 10652 1828
rect 11152 1708 11204 1760
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 1216 1504 1268 1556
rect 11796 1547 11848 1556
rect 11796 1513 11805 1547
rect 11805 1513 11839 1547
rect 11839 1513 11848 1547
rect 11796 1504 11848 1513
rect 13636 1504 13688 1556
rect 16672 1504 16724 1556
rect 11704 1436 11756 1488
rect 13084 1436 13136 1488
rect 18604 1504 18656 1556
rect 3884 1368 3936 1420
rect 11060 1368 11112 1420
rect 3976 1343 4028 1352
rect 3976 1309 3985 1343
rect 3985 1309 4019 1343
rect 4019 1309 4028 1343
rect 3976 1300 4028 1309
rect 13820 1368 13872 1420
rect 14280 1368 14332 1420
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 13820 960 13872 1012
rect 13912 799 13964 808
rect 13912 765 13946 799
rect 13946 765 13964 799
rect 13912 756 13964 765
rect 16120 620 16172 672
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 846 19600 902 20000
rect 2502 19600 2558 20000
rect 4158 19600 4214 20000
rect 5814 19600 5870 20000
rect 7470 19600 7526 20000
rect 9126 19600 9182 20000
rect 10782 19600 10838 20000
rect 12438 19600 12494 20000
rect 14094 19600 14150 20000
rect 15750 19600 15806 20000
rect 17406 19600 17462 20000
rect 19062 19600 19118 20000
rect 860 18834 888 19600
rect 2516 18834 2544 19600
rect 4172 18834 4200 19600
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 5828 18834 5856 19600
rect 7484 18834 7512 19600
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 848 18828 900 18834
rect 848 18770 900 18776
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 2755 18459 3063 18468
rect 4252 18148 4304 18154
rect 4252 18090 4304 18096
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 4264 17882 4292 18090
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4724 17542 4752 18090
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 4804 17808 4856 17814
rect 4804 17750 4856 17756
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 4816 17134 4844 17750
rect 5460 17678 5488 18090
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 4804 17128 4856 17134
rect 4804 17070 4856 17076
rect 2320 16652 2372 16658
rect 2320 16594 2372 16600
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 2332 15570 2360 16594
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 4356 16250 4384 16594
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4816 15910 4844 17070
rect 5460 17066 5488 17614
rect 5644 17610 5672 18090
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 5000 16182 5028 16934
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 5552 16658 5580 17478
rect 5644 16998 5672 17546
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5172 16448 5224 16454
rect 5172 16390 5224 16396
rect 5184 16250 5212 16390
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 4804 15904 4856 15910
rect 4632 15852 4804 15858
rect 4632 15846 4856 15852
rect 4632 15830 4844 15846
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 2332 14550 2360 15506
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 3344 15162 3372 15506
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 3424 15428 3476 15434
rect 3424 15370 3476 15376
rect 3332 15156 3384 15162
rect 3332 15098 3384 15104
rect 3436 14958 3464 15370
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 4264 14618 4292 15438
rect 4356 15366 4384 15506
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 2320 14544 2372 14550
rect 2320 14486 2372 14492
rect 3424 14544 3476 14550
rect 3424 14486 3476 14492
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2148 14074 2176 14418
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2332 12850 2360 14486
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 3252 13870 3280 14418
rect 3436 13870 3464 14486
rect 3620 14006 3648 14554
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3608 14000 3660 14006
rect 3608 13942 3660 13948
rect 3804 13938 3832 14214
rect 4356 13938 4384 15302
rect 4632 14958 4660 15830
rect 5000 15638 5028 16118
rect 5552 15978 5580 16594
rect 5736 16590 5764 17274
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 15978 5764 16526
rect 5540 15972 5592 15978
rect 5540 15914 5592 15920
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 5920 15706 5948 18566
rect 6092 18148 6144 18154
rect 6196 18136 6224 18566
rect 6144 18108 6224 18136
rect 6276 18148 6328 18154
rect 6092 18090 6144 18096
rect 6276 18090 6328 18096
rect 6288 16658 6316 18090
rect 6380 17882 6408 18770
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17882 7420 18226
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 17270 7052 17682
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7392 17066 7420 17478
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 7852 17270 7880 17750
rect 7840 17264 7892 17270
rect 7892 17212 7972 17218
rect 7840 17206 7972 17212
rect 7852 17190 7972 17206
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7392 16794 7420 17002
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6552 16652 6604 16658
rect 6552 16594 6604 16600
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 6012 15638 6040 16186
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6012 15450 6040 15574
rect 6012 15422 6132 15450
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4632 14550 4660 14894
rect 4724 14618 4752 14894
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4620 14544 4672 14550
rect 4620 14486 4672 14492
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4448 14074 4476 14350
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 3792 13932 3844 13938
rect 3792 13874 3844 13880
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3252 13530 3280 13806
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 4172 13326 4200 13806
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2332 12306 2360 12786
rect 2516 12306 2544 13126
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 3804 11218 3832 12786
rect 4172 12442 4200 13262
rect 4632 13190 4660 14486
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5448 14000 5500 14006
rect 5448 13942 5500 13948
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 13394 5028 13670
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 5460 13394 5488 13942
rect 5920 13802 5948 14418
rect 6012 14278 6040 15302
rect 6104 15162 6132 15422
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6288 15026 6316 16594
rect 6564 16250 6592 16594
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 7852 16250 7880 16390
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 16046 7972 17190
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 6380 14482 6408 15846
rect 8036 15434 8064 18566
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8128 17338 8156 17682
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8128 16726 8156 17070
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8128 15570 8156 16458
rect 8220 15978 8248 18022
rect 8208 15972 8260 15978
rect 8208 15914 8260 15920
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 15428 8076 15434
rect 8024 15370 8076 15376
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5552 13530 5580 13738
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4632 12782 4660 13126
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4264 12442 4292 12650
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4252 12436 4304 12442
rect 4252 12378 4304 12384
rect 4816 12306 4844 13126
rect 5460 12986 5488 13330
rect 5920 13326 5948 13738
rect 6196 13394 6224 13806
rect 6472 13462 6500 14418
rect 6656 13870 6684 15098
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 5920 13190 5948 13262
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 6196 12782 6224 13330
rect 6564 13190 6592 13670
rect 6748 13462 6776 14962
rect 7392 14958 7420 15302
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 14074 7328 14350
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7392 13870 7420 14758
rect 8128 14482 8156 15506
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8220 14550 8248 14758
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8404 14482 8432 18838
rect 9140 18834 9168 19600
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8496 17882 8524 18090
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 9600 17626 9628 18022
rect 9692 17746 9720 18294
rect 10152 18222 10180 18634
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 18222 10364 18566
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 18080 10284 18086
rect 10230 18048 10232 18057
rect 10284 18048 10286 18057
rect 9827 17980 10135 17989
rect 10230 17983 10286 17992
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 10336 17678 10364 18158
rect 10324 17672 10376 17678
rect 9600 17598 9720 17626
rect 10324 17614 10376 17620
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8496 16590 8524 16934
rect 9140 16590 9168 16934
rect 9232 16658 9260 17478
rect 9692 17270 9720 17598
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9692 16794 9720 17206
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 10244 16658 10272 17138
rect 10428 17082 10456 18634
rect 10336 17054 10456 17082
rect 10336 16658 10364 17054
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 16726 10456 16934
rect 10416 16720 10468 16726
rect 10416 16662 10468 16668
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 9128 16584 9180 16590
rect 9180 16532 9260 16538
rect 9128 16526 9260 16532
rect 9140 16510 9260 16526
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8496 16114 8524 16390
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 8680 15910 8708 16050
rect 8668 15904 8720 15910
rect 8668 15846 8720 15852
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8496 14482 8524 15642
rect 9048 15570 9076 16050
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9140 15570 9168 15846
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 9232 15502 9260 16510
rect 9496 16516 9548 16522
rect 9496 16458 9548 16464
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9508 16114 9536 16458
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9324 15570 9352 15982
rect 9416 15910 9444 15982
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9600 15570 9628 16050
rect 9692 16046 9720 16458
rect 9876 16250 9904 16594
rect 9968 16454 9996 16594
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9692 15450 9720 15846
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 10244 15706 10272 16594
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10244 15570 10272 15642
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 8588 14958 8616 15438
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8484 14476 8536 14482
rect 8484 14418 8536 14424
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7944 14074 7972 14418
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8036 14074 8064 14350
rect 7932 14068 7984 14074
rect 7932 14010 7984 14016
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8680 14006 8708 15438
rect 9692 15422 9812 15450
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 7380 13864 7432 13870
rect 8300 13864 8352 13870
rect 7380 13806 7432 13812
rect 8220 13824 8300 13852
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13530 6960 13670
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6736 13456 6788 13462
rect 6736 13398 6788 13404
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6184 12776 6236 12782
rect 6104 12736 6184 12764
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 5828 12434 5856 12582
rect 5828 12406 5948 12434
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5736 11898 5764 12242
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5920 11694 5948 12406
rect 6104 11898 6132 12736
rect 6184 12718 6236 12724
rect 6656 12646 6684 13398
rect 6748 12850 6776 13398
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6092 11892 6144 11898
rect 6092 11834 6144 11840
rect 6196 11694 6224 12582
rect 6748 12102 6776 12786
rect 6932 12782 6960 13466
rect 7116 13394 7144 13738
rect 8220 13394 8248 13824
rect 8300 13806 8352 13812
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6932 12442 6960 12718
rect 6920 12436 6972 12442
rect 6920 12378 6972 12384
rect 7116 12306 7144 13194
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 8220 12986 8248 13330
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 7300 12442 7328 12650
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 3988 10810 4016 11154
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3804 10266 3832 10678
rect 5000 10674 5028 10746
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3988 10266 4016 10542
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3884 9920 3936 9926
rect 4264 9897 4292 10066
rect 3884 9862 3936 9868
rect 4250 9888 4306 9897
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 3804 8430 3832 9862
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 3436 7546 3464 7890
rect 3804 7886 3832 8366
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 3620 6458 3648 7278
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3804 6322 3832 7822
rect 3896 7342 3924 9862
rect 4250 9823 4306 9832
rect 4356 9450 4384 10066
rect 4448 9994 4476 10066
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4540 9722 4568 10610
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4632 8634 4660 10542
rect 5460 10470 5488 11562
rect 6840 11354 6868 12106
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6932 10810 6960 11562
rect 8496 11218 8524 13806
rect 8956 13802 8984 14282
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 9232 13394 9260 14214
rect 9416 14074 9444 14350
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9692 13512 9720 15302
rect 9784 14822 9812 15422
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 9692 13484 9812 13512
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9784 13326 9812 13484
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9772 13320 9824 13326
rect 9494 13288 9550 13297
rect 9772 13262 9824 13268
rect 9494 13223 9550 13232
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 8772 10810 8800 11154
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 6184 10736 6236 10742
rect 8484 10736 8536 10742
rect 6236 10696 6500 10724
rect 6184 10678 6236 10684
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9586 4752 9862
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 3976 7948 4028 7954
rect 3976 7890 4028 7896
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3988 5574 4016 7890
rect 4080 7750 4108 8502
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 6662 4108 7686
rect 4172 7342 4200 8230
rect 4264 8090 4292 8366
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4540 7954 4568 8434
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 4724 8294 4752 8366
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4356 7546 4384 7686
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4250 6760 4306 6769
rect 4724 6730 4752 7890
rect 4816 7886 4844 10406
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5092 9586 5120 9930
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5368 9364 5396 10066
rect 5552 9994 5580 10542
rect 6368 10532 6420 10538
rect 6368 10474 6420 10480
rect 6184 10056 6236 10062
rect 5630 10024 5686 10033
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5540 9988 5592 9994
rect 6184 9998 6236 10004
rect 5630 9959 5686 9968
rect 5540 9930 5592 9936
rect 5460 9654 5488 9930
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5368 9336 5488 9364
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 5460 8838 5488 9336
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 5000 8090 5028 8434
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 4988 8084 5040 8090
rect 5040 8044 5120 8072
rect 4988 8026 5040 8032
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7342 4844 7822
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4816 7002 4844 7278
rect 4804 6996 4856 7002
rect 5000 6984 5028 7890
rect 5092 7546 5120 8044
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 4804 6938 4856 6944
rect 4908 6956 5028 6984
rect 5356 6996 5408 7002
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4250 6695 4306 6704
rect 4712 6724 4764 6730
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 5778 4108 6598
rect 4264 5914 4292 6695
rect 4712 6666 4764 6672
rect 4816 6254 4844 6802
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4908 5778 4936 6956
rect 5356 6938 5408 6944
rect 5368 6866 5396 6938
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5368 6746 5396 6802
rect 5276 6718 5396 6746
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6254 5120 6598
rect 5276 6390 5304 6718
rect 5460 6610 5488 7414
rect 5552 7410 5580 9930
rect 5644 9722 5672 9959
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5828 8634 5856 9454
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5632 8356 5684 8362
rect 5632 8298 5684 8304
rect 5644 7954 5672 8298
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5552 6662 5580 7210
rect 5644 6798 5672 7890
rect 5736 7546 5764 7890
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5920 7478 5948 8774
rect 6012 7834 6040 9318
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6104 7954 6132 8366
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6012 7806 6132 7834
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5920 7342 5948 7414
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5368 6582 5488 6610
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5368 6254 5396 6582
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5460 6254 5488 6394
rect 5736 6322 5764 7278
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6322 5948 6734
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6012 6254 6040 6598
rect 5080 6248 5132 6254
rect 5000 6196 5080 6202
rect 5000 6190 5132 6196
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5000 6174 5120 6190
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4908 5574 4936 5714
rect 5000 5710 5028 6174
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 5460 5778 5488 6190
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5816 6112 5868 6118
rect 6104 6066 6132 7806
rect 6196 7546 6224 9998
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6288 9382 6316 9862
rect 6380 9722 6408 10474
rect 6472 9722 6500 10696
rect 8484 10678 8536 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6472 8430 6500 9658
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 9382 6592 9522
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8430 6592 8978
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6288 8294 6316 8366
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6196 6186 6224 7482
rect 6288 7002 6316 7890
rect 6380 7002 6408 8026
rect 6656 7750 6684 10542
rect 6748 10266 6776 10542
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 7024 10062 7052 10406
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6918 9888 6974 9897
rect 6840 9674 6868 9862
rect 6918 9823 6974 9832
rect 6748 9646 6868 9674
rect 6932 9654 6960 9823
rect 6920 9648 6972 9654
rect 6748 9586 6776 9646
rect 6920 9590 6972 9596
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9110 6868 9454
rect 7024 9382 7052 9522
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7116 9178 7144 10542
rect 7208 9722 7236 10542
rect 7484 10266 7512 10542
rect 7668 10266 7696 10610
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 6828 9104 6880 9110
rect 7288 9104 7340 9110
rect 6828 9046 6880 9052
rect 6918 9072 6974 9081
rect 7288 9046 7340 9052
rect 6918 9007 6974 9016
rect 6932 8838 6960 9007
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6748 7954 6776 8434
rect 7012 8424 7064 8430
rect 7012 8366 7064 8372
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6472 7206 6500 7482
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 5816 6054 5868 6060
rect 5552 5846 5580 6054
rect 5644 5914 5672 6054
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5828 5778 5856 6054
rect 6012 6038 6132 6066
rect 6012 5778 6040 6038
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 3988 4078 4016 5510
rect 5092 5302 5120 5714
rect 5828 5658 5856 5714
rect 5552 5630 5856 5658
rect 5552 5574 5580 5630
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5828 5030 5856 5510
rect 6012 5098 6040 5714
rect 6196 5710 6224 6122
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 3700 2916 3752 2922
rect 3700 2858 3752 2864
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 1216 1556 1268 1562
rect 1216 1498 1268 1504
rect 1228 400 1256 1498
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 3712 400 3740 2858
rect 3882 1456 3938 1465
rect 3882 1391 3884 1400
rect 3936 1391 3938 1400
rect 3884 1362 3936 1368
rect 3988 1358 4016 4014
rect 5644 4010 5672 4966
rect 6380 4690 6408 6938
rect 6748 6322 6776 7414
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6472 5370 6500 5510
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6564 5234 6592 5510
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6656 5098 6684 5306
rect 6840 5273 6868 5714
rect 6826 5264 6882 5273
rect 6826 5199 6882 5208
rect 6932 5166 6960 7890
rect 7024 6866 7052 8366
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7116 7342 7144 8230
rect 7208 8090 7236 8366
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7116 6458 7144 7142
rect 7208 6866 7236 7210
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7208 6304 7236 6802
rect 7300 6798 7328 9046
rect 7392 8838 7420 10202
rect 8036 9994 8064 10406
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 8036 9586 8064 9930
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7562 9208 7618 9217
rect 7668 9178 7696 9454
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 7562 9143 7618 9152
rect 7656 9172 7708 9178
rect 7576 9042 7604 9143
rect 7656 9114 7708 9120
rect 7760 9110 7788 9318
rect 7748 9104 7800 9110
rect 7748 9046 7800 9052
rect 7930 9072 7986 9081
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7840 9036 7892 9042
rect 8036 9058 8064 9522
rect 8128 9178 8156 10066
rect 8220 10033 8248 10066
rect 8206 10024 8262 10033
rect 8206 9959 8262 9968
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 8036 9030 8156 9058
rect 7930 9007 7986 9016
rect 7840 8978 7892 8984
rect 7852 8945 7880 8978
rect 7838 8936 7894 8945
rect 7944 8906 7972 9007
rect 7838 8871 7894 8880
rect 7932 8900 7984 8906
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 7852 8498 7880 8871
rect 7932 8842 7984 8848
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7944 7750 7972 8366
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7484 6905 7512 7414
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7470 6896 7526 6905
rect 7668 6866 7696 7142
rect 7470 6831 7472 6840
rect 7524 6831 7526 6840
rect 7656 6860 7708 6866
rect 7472 6802 7524 6808
rect 7656 6802 7708 6808
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7116 6276 7236 6304
rect 7116 5574 7144 6276
rect 7300 6202 7328 6734
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6254 7420 6598
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 7852 6254 7880 7414
rect 7944 7410 7972 7686
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8036 7290 8064 8774
rect 7944 7262 8064 7290
rect 7944 6730 7972 7262
rect 8128 6746 8156 9030
rect 8220 8838 8248 9590
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 7342 8248 8774
rect 8312 8294 8340 10202
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 7410 8340 8230
rect 8404 7546 8432 10134
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 6934 8248 7278
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8208 6792 8260 6798
rect 8128 6740 8208 6746
rect 8128 6734 8260 6740
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 8024 6724 8076 6730
rect 8128 6718 8248 6734
rect 8024 6666 8076 6672
rect 7944 6254 7972 6666
rect 7208 6174 7328 6202
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7208 5778 7236 6174
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7300 5166 7328 6054
rect 7392 5778 7420 6190
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 5658 7604 5714
rect 7852 5710 7880 6190
rect 8036 6118 8064 6666
rect 8220 6458 8248 6718
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8220 6186 8248 6394
rect 8312 6390 8340 7346
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7392 5642 7604 5658
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 7380 5636 7604 5642
rect 7432 5630 7604 5636
rect 7380 5578 7432 5584
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6644 5092 6696 5098
rect 6644 5034 6696 5040
rect 6932 4826 6960 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7392 4758 7420 5578
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7380 4752 7432 4758
rect 7380 4694 7432 4700
rect 7760 4690 7788 5102
rect 7852 4826 7880 5646
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7944 4690 7972 4966
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7472 4616 7524 4622
rect 7392 4564 7472 4570
rect 7392 4558 7524 4564
rect 7852 4570 7880 4626
rect 8036 4570 8064 4966
rect 7392 4542 7512 4558
rect 7852 4542 8064 4570
rect 7392 4214 7420 4542
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 7380 4208 7432 4214
rect 8220 4185 8248 4422
rect 7380 4150 7432 4156
rect 8206 4176 8262 4185
rect 8206 4111 8262 4120
rect 8312 4078 8340 5646
rect 8404 4690 8432 7482
rect 8496 7274 8524 10678
rect 8772 10062 8800 10746
rect 9416 10606 9444 12922
rect 9508 12714 9536 13223
rect 9876 13002 9904 13398
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9692 12974 9904 13002
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9508 11082 9536 11630
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 10810 9536 11018
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9416 10130 9444 10542
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 9416 9586 9444 10066
rect 9692 9654 9720 12974
rect 9772 12912 9824 12918
rect 9770 12880 9772 12889
rect 9824 12880 9826 12889
rect 9770 12815 9826 12824
rect 9968 12782 9996 13330
rect 10048 13320 10100 13326
rect 10244 13274 10272 14758
rect 10336 14482 10364 16594
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10428 15638 10456 15846
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10520 15570 10548 18906
rect 10796 18834 10824 19600
rect 12452 18834 12480 19600
rect 14108 18834 14136 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 15764 18834 15792 19600
rect 17420 18834 17448 19600
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10612 17202 10640 17818
rect 10796 17678 10824 18294
rect 11060 18148 11112 18154
rect 11060 18090 11112 18096
rect 11072 17882 11100 18090
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11900 17746 11928 18362
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10612 13326 10640 16730
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10704 16454 10732 16662
rect 10980 16454 11008 17070
rect 11072 17066 11100 17546
rect 11612 17196 11664 17202
rect 11612 17138 11664 17144
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11072 16522 11100 17002
rect 11060 16516 11112 16522
rect 11060 16458 11112 16464
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16182 11008 16390
rect 11072 16182 11100 16458
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10980 15706 11008 15982
rect 10968 15700 11020 15706
rect 10968 15642 11020 15648
rect 11072 14618 11100 16118
rect 11624 16046 11652 17138
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11520 15972 11572 15978
rect 11520 15914 11572 15920
rect 11532 15706 11560 15914
rect 11520 15700 11572 15706
rect 11520 15642 11572 15648
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 14958 11284 15506
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10048 13262 10100 13268
rect 10060 13161 10088 13262
rect 10152 13246 10272 13274
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10690 13288 10746 13297
rect 10046 13152 10102 13161
rect 10046 13087 10102 13096
rect 10060 12782 10088 13087
rect 10152 13025 10180 13246
rect 10690 13223 10746 13232
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10138 13016 10194 13025
rect 10138 12951 10140 12960
rect 10192 12951 10194 12960
rect 10140 12922 10192 12928
rect 10244 12782 10272 13126
rect 10704 12918 10732 13223
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 9956 12776 10008 12782
rect 9954 12744 9956 12753
rect 10048 12776 10100 12782
rect 10008 12744 10010 12753
rect 10048 12718 10100 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 9954 12679 10010 12688
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10470 9904 10950
rect 10060 10674 10088 11290
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8588 9110 8616 9318
rect 8758 9208 8814 9217
rect 8758 9143 8814 9152
rect 8576 9104 8628 9110
rect 8668 9104 8720 9110
rect 8576 9046 8628 9052
rect 8666 9072 8668 9081
rect 8720 9072 8722 9081
rect 8772 9042 8800 9143
rect 8666 9007 8722 9016
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8668 8968 8720 8974
rect 8666 8936 8668 8945
rect 8944 8968 8996 8974
rect 8720 8936 8722 8945
rect 8944 8910 8996 8916
rect 8666 8871 8722 8880
rect 8956 8362 8984 8910
rect 9048 8838 9076 9318
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9140 8634 9168 9046
rect 9232 8974 9260 9454
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 9042 9536 9386
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9508 8634 9536 8978
rect 9600 8945 9628 8978
rect 9586 8936 9642 8945
rect 9586 8871 9642 8880
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9508 8022 9536 8298
rect 9600 8090 9628 8366
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 8484 7268 8536 7274
rect 8484 7210 8536 7216
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 8666 6896 8722 6905
rect 8666 6831 8668 6840
rect 8720 6831 8722 6840
rect 8668 6802 8720 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6322 8524 6598
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 8496 5302 8524 6054
rect 8588 5710 8616 6734
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8484 5296 8536 5302
rect 8576 5296 8628 5302
rect 8484 5238 8536 5244
rect 8574 5264 8576 5273
rect 8628 5264 8630 5273
rect 8496 5166 8524 5238
rect 8680 5234 8708 6802
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8574 5199 8630 5208
rect 8668 5228 8720 5234
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8496 4570 8524 5102
rect 8588 4758 8616 5199
rect 8668 5170 8720 5176
rect 8956 5166 8984 6394
rect 9324 5778 9352 7210
rect 9692 6254 9720 9590
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8838 9812 8978
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9968 8566 9996 8842
rect 10152 8634 10180 9114
rect 10244 9058 10272 12038
rect 10336 11830 10364 12854
rect 10506 12744 10562 12753
rect 10796 12730 10824 14214
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 11058 13152 11114 13161
rect 10874 13016 10930 13025
rect 10874 12951 10930 12960
rect 10506 12679 10562 12688
rect 10612 12702 10824 12730
rect 10416 12640 10468 12646
rect 10414 12608 10416 12617
rect 10468 12608 10470 12617
rect 10414 12543 10470 12552
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 11354 10364 11630
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 9178 10364 10950
rect 10428 10606 10456 12543
rect 10416 10600 10468 10606
rect 10416 10542 10468 10548
rect 10520 10538 10548 12679
rect 10612 12646 10640 12702
rect 10600 12640 10652 12646
rect 10784 12640 10836 12646
rect 10600 12582 10652 12588
rect 10782 12608 10784 12617
rect 10836 12608 10838 12617
rect 10782 12543 10838 12552
rect 10784 12368 10836 12374
rect 10782 12336 10784 12345
rect 10836 12336 10838 12345
rect 10600 12300 10652 12306
rect 10782 12271 10838 12280
rect 10600 12242 10652 12248
rect 10612 11898 10640 12242
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10520 9674 10548 10474
rect 10428 9646 10548 9674
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10244 9030 10364 9058
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 10046 8528 10102 8537
rect 9784 8401 9812 8502
rect 10152 8498 10180 8570
rect 10046 8463 10102 8472
rect 10140 8492 10192 8498
rect 9956 8424 10008 8430
rect 9770 8392 9826 8401
rect 9770 8327 9826 8336
rect 9954 8392 9956 8401
rect 10008 8392 10010 8401
rect 9954 8327 10010 8336
rect 10060 8294 10088 8463
rect 10140 8434 10192 8440
rect 10244 8362 10272 8910
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9770 7984 9826 7993
rect 10152 7954 10180 8026
rect 9770 7919 9772 7928
rect 9824 7919 9826 7928
rect 10140 7948 10192 7954
rect 9772 7890 9824 7896
rect 10140 7890 10192 7896
rect 10244 7818 10272 8298
rect 10232 7812 10284 7818
rect 10232 7754 10284 7760
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9416 5710 9444 6054
rect 9692 5914 9720 6190
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9404 5568 9456 5574
rect 9508 5556 9536 5714
rect 9456 5528 9536 5556
rect 9404 5510 9456 5516
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8496 4542 8616 4570
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4078 8432 4422
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 7208 3670 7236 3878
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 8312 3602 8340 4014
rect 8588 3602 8616 4542
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4282 8708 4422
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8956 4214 8984 5102
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8956 4010 8984 4150
rect 8944 4004 8996 4010
rect 8944 3946 8996 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3602 9720 3878
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 6196 400 6224 2790
rect 10336 2774 10364 9030
rect 10428 8906 10456 9646
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10520 8566 10548 9318
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10508 8560 10560 8566
rect 10508 8502 10560 8508
rect 10612 8430 10640 8570
rect 10416 8424 10468 8430
rect 10600 8424 10652 8430
rect 10468 8401 10548 8412
rect 10468 8392 10562 8401
rect 10468 8384 10506 8392
rect 10416 8366 10468 8372
rect 10600 8366 10652 8372
rect 10506 8327 10562 8336
rect 10414 8256 10470 8265
rect 10414 8191 10470 8200
rect 10428 6730 10456 8191
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7342 10548 7686
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10520 6866 10548 7278
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10520 6769 10548 6802
rect 10506 6760 10562 6769
rect 10416 6724 10468 6730
rect 10506 6695 10562 6704
rect 10416 6666 10468 6672
rect 10704 2774 10732 11766
rect 10888 11354 10916 12951
rect 10980 12714 11008 13126
rect 11058 13087 11114 13096
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10980 12374 11008 12650
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10606 10824 11154
rect 10888 11014 10916 11290
rect 10980 11121 11008 12038
rect 11072 11218 11100 13087
rect 11164 12442 11192 14826
rect 11348 14482 11376 15370
rect 11808 14958 11836 15982
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 11256 13802 11284 14418
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11348 13841 11376 13942
rect 11334 13832 11390 13841
rect 11244 13796 11296 13802
rect 11334 13767 11390 13776
rect 11244 13738 11296 13744
rect 11152 12436 11204 12442
rect 11440 12434 11468 13942
rect 11532 13802 11560 14214
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11532 12442 11560 12922
rect 11152 12378 11204 12384
rect 11348 12406 11468 12434
rect 11520 12436 11572 12442
rect 11244 11280 11296 11286
rect 11244 11222 11296 11228
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10966 11112 11022 11121
rect 10966 11047 11022 11056
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10606 10916 10950
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10796 8537 10824 10542
rect 11256 10470 11284 11222
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10888 8566 10916 9386
rect 10980 9382 11008 10406
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9722 11192 10066
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11058 9616 11114 9625
rect 11058 9551 11114 9560
rect 11072 9518 11100 9551
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10980 8566 11008 8978
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10876 8560 10928 8566
rect 10782 8528 10838 8537
rect 10876 8502 10928 8508
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 11072 8514 11100 8842
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10782 8463 10838 8472
rect 10796 8294 10824 8463
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10980 8090 11008 8502
rect 11072 8486 11192 8514
rect 11058 8392 11114 8401
rect 11058 8327 11060 8336
rect 11112 8327 11114 8336
rect 11060 8298 11112 8304
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10888 6934 10916 7958
rect 11072 7002 11100 8298
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10888 5234 10916 6870
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4690 10916 5170
rect 10980 4826 11008 6938
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11072 5098 11100 5306
rect 11164 5302 11192 8486
rect 11256 6662 11284 8774
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6186 11284 6598
rect 11244 6180 11296 6186
rect 11244 6122 11296 6128
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11256 5166 11284 6122
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 3738 10916 4626
rect 11150 4176 11206 4185
rect 11150 4111 11206 4120
rect 11164 4010 11192 4111
rect 11348 4010 11376 12406
rect 11624 12434 11652 12922
rect 11716 12646 11744 14758
rect 11992 12918 12020 18566
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12084 16454 12112 18158
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12256 17196 12308 17202
rect 12256 17138 12308 17144
rect 12268 16658 12296 17138
rect 12360 16726 12388 17274
rect 12348 16720 12400 16726
rect 12348 16662 12400 16668
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16046 12112 16390
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 15366 12112 15982
rect 12544 15978 12572 18634
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 17882 12664 18090
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12820 17746 12848 18566
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12912 17270 12940 17682
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 14414 12112 15302
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 12544 15026 12572 15914
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12544 14482 12572 14962
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 13938 12112 14350
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12084 13530 12112 13874
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11808 12753 11836 12854
rect 11794 12744 11850 12753
rect 11794 12679 11850 12688
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11624 12406 11744 12434
rect 11520 12378 11572 12384
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10130 11468 10950
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11440 9178 11468 10066
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11532 9042 11560 10066
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11624 9518 11652 9590
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11440 8362 11468 8570
rect 11624 8548 11652 9454
rect 11532 8520 11652 8548
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11532 7410 11560 8520
rect 11612 8288 11664 8294
rect 11610 8256 11612 8265
rect 11664 8256 11666 8265
rect 11610 8191 11666 8200
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11428 6724 11480 6730
rect 11428 6666 11480 6672
rect 11440 6390 11468 6666
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11440 4078 11468 5510
rect 11532 5030 11560 7346
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 6458 11652 6802
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4690 11560 4966
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11428 4072 11480 4078
rect 11428 4014 11480 4020
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 11440 3670 11468 4014
rect 11532 3942 11560 4626
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 10244 2746 10364 2774
rect 10612 2746 10732 2774
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 8680 400 8708 2586
rect 10244 2582 10272 2746
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10612 1834 10640 2746
rect 11072 2446 11100 3606
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11072 1902 11100 2382
rect 11060 1896 11112 1902
rect 11060 1838 11112 1844
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 11072 1426 11100 1838
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 11164 400 11192 1702
rect 11716 1494 11744 12406
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11796 11620 11848 11626
rect 11796 11562 11848 11568
rect 11808 11286 11836 11562
rect 11900 11354 11928 12174
rect 12084 11830 12112 13466
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12782 12388 12854
rect 12544 12850 12572 13670
rect 12636 13394 12664 16934
rect 13004 16794 13032 17070
rect 13556 17066 13584 18566
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 15120 17202 15148 17614
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 13556 16046 13584 17002
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 16132 16250 16160 18566
rect 16684 18222 16712 18566
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17134 16620 18022
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13096 15570 13124 15846
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14550 13124 14894
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13734 12848 13806
rect 12808 13728 12860 13734
rect 12808 13670 12860 13676
rect 12820 13530 12848 13670
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12532 12844 12584 12850
rect 12532 12786 12584 12792
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12256 11620 12308 11626
rect 12256 11562 12308 11568
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11900 9217 11928 10406
rect 12084 10266 12112 11154
rect 12268 11014 12296 11562
rect 12452 11098 12480 11698
rect 12544 11558 12572 12242
rect 12636 11694 12664 12310
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12728 11121 12756 12174
rect 12714 11112 12770 11121
rect 12452 11070 12572 11098
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 9722 12112 9998
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12452 9602 12480 9658
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12360 9574 12480 9602
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11886 9208 11942 9217
rect 11886 9143 11942 9152
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 6662 11928 8366
rect 11992 8090 12020 8978
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11992 7546 12020 8026
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11992 7206 12020 7482
rect 12084 7274 12112 9386
rect 12268 8945 12296 9522
rect 12360 9518 12388 9574
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12452 9382 12480 9454
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 8974 12480 9318
rect 12440 8968 12492 8974
rect 12254 8936 12310 8945
rect 12440 8910 12492 8916
rect 12254 8871 12310 8880
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 12254 7440 12310 7449
rect 12254 7375 12310 7384
rect 12268 7342 12296 7375
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 12084 6984 12112 7210
rect 12176 7002 12204 7278
rect 11992 6956 12112 6984
rect 12164 6996 12216 7002
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6254 11928 6598
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11808 6118 11836 6190
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11900 5642 11928 6190
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 11992 5370 12020 6956
rect 12164 6938 12216 6944
rect 12268 6866 12296 7278
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12084 6390 12112 6802
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 4865 12020 5306
rect 12084 5234 12112 6326
rect 12544 5914 12572 11070
rect 12714 11047 12770 11056
rect 12716 10192 12768 10198
rect 12716 10134 12768 10140
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12636 9042 12664 9522
rect 12728 9489 12756 10134
rect 12808 9512 12860 9518
rect 12714 9480 12770 9489
rect 12808 9454 12860 9460
rect 12912 9466 12940 13874
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 12306 13032 13670
rect 13096 12782 13124 14486
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13372 13870 13400 14418
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13188 12889 13216 13330
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13188 11694 13216 12815
rect 13464 11898 13492 13874
rect 13556 12714 13584 15846
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13648 14006 13676 14554
rect 13832 14074 13860 14894
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13924 14482 13952 14758
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13648 13818 13676 13942
rect 13648 13790 13768 13818
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13648 13394 13676 13670
rect 13740 13394 13768 13790
rect 13924 13394 13952 14214
rect 14016 13938 14044 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 14476 13530 14504 14010
rect 14936 13870 14964 14282
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13728 13388 13780 13394
rect 13728 13330 13780 13336
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13832 12442 13860 12718
rect 14476 12442 14504 13466
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13452 11892 13504 11898
rect 13452 11834 13504 11840
rect 13280 11694 13308 11834
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13464 11626 13492 11834
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 9586 13032 10406
rect 13188 10130 13216 10610
rect 13464 10266 13492 11154
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12714 9415 12770 9424
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12728 9178 12756 9318
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8566 12664 8774
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12820 8022 12848 9454
rect 12912 9438 13032 9466
rect 13004 9058 13032 9438
rect 13096 9382 13124 10066
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9722 13216 9862
rect 13280 9722 13308 9998
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13464 9654 13492 10066
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13266 9208 13322 9217
rect 13266 9143 13322 9152
rect 12912 9030 13032 9058
rect 13174 9072 13230 9081
rect 13280 9042 13308 9143
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12636 6866 12664 7754
rect 12728 7002 12756 7822
rect 12912 7546 12940 9030
rect 13174 9007 13176 9016
rect 13228 9007 13230 9016
rect 13268 9036 13320 9042
rect 13176 8978 13228 8984
rect 13268 8978 13320 8984
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 12992 8968 13044 8974
rect 12990 8936 12992 8945
rect 13044 8936 13046 8945
rect 12990 8871 13046 8880
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12820 6866 12848 7414
rect 13004 7410 13032 8871
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13096 7886 13124 8774
rect 13084 7880 13136 7886
rect 13084 7822 13136 7828
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12912 7002 12940 7278
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 13096 6118 13124 7822
rect 13188 6322 13216 8978
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13280 7342 13308 8434
rect 13372 8090 13400 8910
rect 13464 8566 13492 8978
rect 13556 8634 13584 12174
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13740 11354 13768 11562
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13832 11218 13860 12106
rect 14016 11354 14044 12106
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 14292 11150 14320 11630
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11218 14412 11494
rect 14476 11354 14504 11562
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13912 10056 13964 10062
rect 13740 10004 13912 10010
rect 13740 9998 13964 10004
rect 13740 9982 13952 9998
rect 13740 9926 13768 9982
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13728 9512 13780 9518
rect 13832 9500 13860 9862
rect 14016 9518 14044 9862
rect 13780 9472 13860 9500
rect 14004 9512 14056 9518
rect 13728 9454 13780 9460
rect 14004 9454 14056 9460
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 8974 13676 9318
rect 13740 9042 13768 9454
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13832 8838 13860 9318
rect 14016 9217 14044 9318
rect 14002 9208 14058 9217
rect 14002 9143 14058 9152
rect 14108 9042 14136 10066
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 9178 14228 9454
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14292 9058 14320 11086
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 14832 10124 14884 10130
rect 14832 10066 14884 10072
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14384 9450 14412 9998
rect 14844 9722 14872 10066
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 9444 14424 9450
rect 14372 9386 14424 9392
rect 14384 9178 14412 9386
rect 14372 9172 14424 9178
rect 14372 9114 14424 9120
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14200 9030 14320 9058
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 13924 8090 13952 8298
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 7528 13584 7822
rect 13636 7540 13688 7546
rect 13556 7500 13636 7528
rect 13268 7336 13320 7342
rect 13268 7278 13320 7284
rect 13280 6866 13308 7278
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13464 6662 13492 7210
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 13464 5778 13492 6598
rect 13556 6254 13584 7500
rect 13636 7482 13688 7488
rect 13832 7342 13860 7890
rect 14016 7750 14044 8298
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14108 7449 14136 8978
rect 14200 8430 14228 9030
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14292 8566 14320 8774
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14094 7440 14150 7449
rect 14094 7375 14150 7384
rect 13820 7336 13872 7342
rect 14200 7324 14228 8366
rect 13820 7278 13872 7284
rect 14108 7296 14228 7324
rect 13832 6866 13860 7278
rect 13820 6860 13872 6866
rect 13872 6820 13952 6848
rect 13820 6802 13872 6808
rect 13924 6254 13952 6820
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 12898 5400 12954 5409
rect 12898 5335 12900 5344
rect 12952 5335 12954 5344
rect 12900 5306 12952 5312
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 11978 4856 12034 4865
rect 12452 4826 12480 5102
rect 12728 4826 12756 5102
rect 11978 4791 12034 4800
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12360 4706 12388 4762
rect 11980 4684 12032 4690
rect 12360 4678 12480 4706
rect 11980 4626 12032 4632
rect 11992 4282 12020 4626
rect 12452 4622 12480 4678
rect 12716 4684 12768 4690
rect 12820 4672 12848 5238
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4826 12940 4966
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12768 4644 12848 4672
rect 12716 4626 12768 4632
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12728 4554 12756 4626
rect 12716 4548 12768 4554
rect 12716 4490 12768 4496
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12912 4282 12940 4422
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12820 3738 12848 4014
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 13004 3398 13032 5714
rect 13096 5030 13124 5714
rect 13188 5370 13216 5714
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 13096 4758 13124 4966
rect 13174 4856 13230 4865
rect 13280 4842 13308 5646
rect 13556 5137 13584 6190
rect 13832 6118 13860 6190
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5642 13860 6054
rect 14108 5914 14136 7296
rect 14292 6254 14320 8366
rect 14384 7818 14412 9114
rect 14476 8906 14504 9454
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14936 9042 14964 11494
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 14924 9036 14976 9042
rect 14924 8978 14976 8984
rect 15028 8974 15056 10542
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14280 6248 14332 6254
rect 14332 6196 14412 6202
rect 14280 6190 14412 6196
rect 14292 6174 14412 6190
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14002 5808 14058 5817
rect 14002 5743 14004 5752
rect 14056 5743 14058 5752
rect 14004 5714 14056 5720
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 14200 5166 14228 6054
rect 14292 5846 14320 6054
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14384 5386 14412 6174
rect 14476 5778 14504 8298
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6390 14688 6598
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 14936 5914 14964 8570
rect 15028 7954 15056 8910
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15016 6180 15068 6186
rect 15016 6122 15068 6128
rect 15028 5914 15056 6122
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15016 5908 15068 5914
rect 15016 5850 15068 5856
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15028 5642 15056 5714
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14292 5358 14412 5386
rect 13820 5160 13872 5166
rect 13542 5128 13598 5137
rect 13820 5102 13872 5108
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13542 5063 13598 5072
rect 13230 4814 13308 4842
rect 13174 4791 13230 4800
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13188 4622 13216 4791
rect 13176 4616 13228 4622
rect 13176 4558 13228 4564
rect 13188 4146 13216 4558
rect 13556 4554 13584 5063
rect 13832 4554 13860 5102
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4690 14136 4966
rect 14096 4684 14148 4690
rect 14200 4672 14228 5102
rect 14292 4826 14320 5358
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 5114 14412 5170
rect 14384 5086 14504 5114
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4820 14332 4826
rect 14280 4762 14332 4768
rect 14280 4684 14332 4690
rect 14200 4644 14280 4672
rect 14096 4626 14148 4632
rect 14280 4626 14332 4632
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14108 4570 14136 4626
rect 14384 4570 14412 4966
rect 14476 4826 14504 5086
rect 14660 5030 14688 5510
rect 14936 5234 14964 5510
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14936 4690 14964 4966
rect 14556 4684 14608 4690
rect 14556 4626 14608 4632
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 13544 4548 13596 4554
rect 13544 4490 13596 4496
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13740 4078 13768 4218
rect 13832 4214 13860 4490
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 14016 4010 14044 4558
rect 14108 4542 14412 4570
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14476 4282 14504 4558
rect 14568 4282 14596 4626
rect 14752 4554 14780 4626
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14936 4146 14964 4626
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15028 4078 15056 4966
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14004 4004 14056 4010
rect 14004 3946 14056 3952
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 11808 1562 11836 2790
rect 12820 2650 12848 2790
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 13082 2680 13138 2689
rect 14542 2683 14850 2692
rect 12808 2644 12860 2650
rect 13082 2615 13138 2624
rect 12808 2586 12860 2592
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 11796 1556 11848 1562
rect 11796 1498 11848 1504
rect 13096 1494 13124 2615
rect 15120 2582 15148 12854
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15304 10674 15608 10690
rect 15292 10668 15608 10674
rect 15344 10662 15608 10668
rect 15292 10610 15344 10616
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9654 15240 10066
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15200 9512 15252 9518
rect 15198 9480 15200 9489
rect 15252 9480 15254 9489
rect 15198 9415 15254 9424
rect 15212 7954 15240 9415
rect 15304 9081 15332 10610
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10130 15424 10542
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15290 9072 15346 9081
rect 15396 9042 15424 9318
rect 15290 9007 15346 9016
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15396 8430 15424 8978
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15488 8294 15516 10134
rect 15580 10130 15608 10662
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15580 9450 15608 9862
rect 15856 9654 15884 11222
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8634 15608 8774
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15200 7948 15252 7954
rect 15384 7948 15436 7954
rect 15252 7908 15332 7936
rect 15200 7890 15252 7896
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 6202 15240 7210
rect 15304 6304 15332 7908
rect 15384 7890 15436 7896
rect 15396 7274 15424 7890
rect 15488 7342 15516 8230
rect 15580 7954 15608 8570
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 6798 15424 7210
rect 15476 6996 15528 7002
rect 15672 6984 15700 9590
rect 16040 9586 16068 10406
rect 16224 10266 16252 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16132 9518 16160 10066
rect 16500 9518 16528 10066
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15948 8974 15976 9318
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 16132 8922 16160 9454
rect 16224 9042 16252 9454
rect 16408 9382 16436 9454
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 15948 8480 15976 8910
rect 16132 8894 16252 8922
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16028 8492 16080 8498
rect 15948 8452 16028 8480
rect 15948 7954 15976 8452
rect 16028 8434 16080 8440
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15764 7546 15792 7890
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15948 7410 15976 7686
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15528 6956 15700 6984
rect 15476 6938 15528 6944
rect 15488 6798 15516 6938
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15488 6338 15516 6734
rect 15580 6458 15608 6734
rect 15672 6458 15700 6802
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15488 6310 15608 6338
rect 15304 6276 15424 6304
rect 15212 6186 15332 6202
rect 15212 6180 15344 6186
rect 15212 6174 15292 6180
rect 15292 6122 15344 6128
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5166 15240 6054
rect 15396 5234 15424 6276
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5710 15516 6190
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15488 5370 15516 5646
rect 15580 5642 15608 6310
rect 15672 5778 15700 6394
rect 15948 6322 15976 6802
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16132 6254 16160 8774
rect 16224 8634 16252 8894
rect 16408 8838 16436 9318
rect 16500 9024 16528 9454
rect 16580 9444 16632 9450
rect 16580 9386 16632 9392
rect 16592 9178 16620 9386
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16580 9036 16632 9042
rect 16500 8996 16580 9024
rect 16580 8978 16632 8984
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16028 6248 16080 6254
rect 16028 6190 16080 6196
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16040 6118 16068 6190
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16026 5808 16082 5817
rect 15660 5772 15712 5778
rect 16026 5743 16028 5752
rect 15660 5714 15712 5720
rect 16080 5743 16082 5752
rect 16028 5714 16080 5720
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15396 4672 15424 5170
rect 15476 5160 15528 5166
rect 15474 5128 15476 5137
rect 15528 5128 15530 5137
rect 15474 5063 15530 5072
rect 15580 4690 15608 5578
rect 16040 5370 16068 5714
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16132 4690 16160 6190
rect 16224 5817 16252 8026
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16316 6458 16344 7890
rect 16408 6866 16436 8298
rect 16592 8022 16620 8842
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16500 7546 16528 7890
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16488 7540 16540 7546
rect 16488 7482 16540 7488
rect 16488 7336 16540 7342
rect 16592 7324 16620 7822
rect 16540 7296 16620 7324
rect 16488 7278 16540 7284
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16302 6352 16358 6361
rect 16408 6322 16436 6802
rect 16500 6361 16528 7278
rect 16486 6352 16542 6361
rect 16302 6287 16358 6296
rect 16396 6316 16448 6322
rect 16210 5808 16266 5817
rect 16210 5743 16266 5752
rect 16212 5636 16264 5642
rect 16212 5578 16264 5584
rect 16224 5166 16252 5578
rect 16316 5166 16344 6287
rect 16486 6287 16542 6296
rect 16396 6258 16448 6264
rect 16408 6202 16436 6258
rect 16408 6174 16528 6202
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5778 16436 6054
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16500 5166 16528 6174
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16592 5778 16620 6122
rect 16580 5772 16632 5778
rect 16580 5714 16632 5720
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 15476 4684 15528 4690
rect 15396 4644 15476 4672
rect 15476 4626 15528 4632
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16316 4214 16344 5102
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 14280 2440 14332 2446
rect 14280 2382 14332 2388
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 11704 1488 11756 1494
rect 11704 1430 11756 1436
rect 13084 1488 13136 1494
rect 13084 1430 13136 1436
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 13648 400 13676 1498
rect 14292 1426 14320 2382
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 16684 1562 16712 13126
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 19076 9625 19104 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 19062 9616 19118 9625
rect 19062 9551 19118 9560
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 8838 16804 9318
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16776 8430 16804 8774
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 17236 8634 17264 8978
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 16764 8424 16816 8430
rect 16764 8366 16816 8372
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16776 7954 16804 8026
rect 17236 8022 17264 8570
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16764 7812 16816 7818
rect 16764 7754 16816 7760
rect 16776 7342 16804 7754
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 17224 6180 17276 6186
rect 17224 6122 17276 6128
rect 17236 5778 17264 6122
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 16672 1556 16724 1562
rect 16672 1498 16724 1504
rect 18604 1556 18656 1562
rect 18604 1498 18656 1504
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14280 1420 14332 1426
rect 14280 1362 14332 1368
rect 13832 1018 13860 1362
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 13820 1012 13872 1018
rect 13820 954 13872 960
rect 13910 912 13966 921
rect 13910 847 13966 856
rect 13924 814 13952 847
rect 13912 808 13964 814
rect 13912 750 13964 756
rect 16120 672 16172 678
rect 16120 614 16172 620
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 16132 400 16160 614
rect 18616 400 18644 1498
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
rect 11150 0 11206 400
rect 13634 0 13690 400
rect 16118 0 16174 400
rect 18602 0 18658 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 10230 18028 10232 18048
rect 10232 18028 10284 18048
rect 10284 18028 10286 18048
rect 10230 17992 10286 18028
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 4250 9832 4306 9888
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 9494 13232 9550 13288
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 4250 6704 4306 6760
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 5630 9968 5686 10024
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 6918 9832 6974 9888
rect 6918 9016 6974 9072
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 3882 1420 3938 1456
rect 3882 1400 3884 1420
rect 3884 1400 3936 1420
rect 3936 1400 3938 1420
rect 6826 5208 6882 5264
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 7562 9152 7618 9208
rect 7930 9016 7986 9072
rect 8206 9968 8262 10024
rect 7838 8880 7894 8936
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 7470 6860 7526 6896
rect 7470 6840 7472 6860
rect 7472 6840 7524 6860
rect 7524 6840 7526 6860
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 8206 4120 8262 4176
rect 9770 12860 9772 12880
rect 9772 12860 9824 12880
rect 9824 12860 9826 12880
rect 9770 12824 9826 12860
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 10046 13096 10102 13152
rect 10690 13232 10746 13288
rect 10138 12980 10194 13016
rect 10138 12960 10140 12980
rect 10140 12960 10192 12980
rect 10192 12960 10194 12980
rect 9954 12724 9956 12744
rect 9956 12724 10008 12744
rect 10008 12724 10010 12744
rect 9954 12688 10010 12724
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 8758 9152 8814 9208
rect 8666 9052 8668 9072
rect 8668 9052 8720 9072
rect 8720 9052 8722 9072
rect 8666 9016 8722 9052
rect 8666 8916 8668 8936
rect 8668 8916 8720 8936
rect 8720 8916 8722 8936
rect 8666 8880 8722 8916
rect 9586 8880 9642 8936
rect 8666 6860 8722 6896
rect 8666 6840 8668 6860
rect 8668 6840 8720 6860
rect 8720 6840 8722 6860
rect 8574 5244 8576 5264
rect 8576 5244 8628 5264
rect 8628 5244 8630 5264
rect 8574 5208 8630 5244
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 10506 12688 10562 12744
rect 10874 12960 10930 13016
rect 10414 12588 10416 12608
rect 10416 12588 10468 12608
rect 10468 12588 10470 12608
rect 10414 12552 10470 12588
rect 10782 12588 10784 12608
rect 10784 12588 10836 12608
rect 10836 12588 10838 12608
rect 10782 12552 10838 12588
rect 10782 12316 10784 12336
rect 10784 12316 10836 12336
rect 10836 12316 10838 12336
rect 10782 12280 10838 12316
rect 10046 8472 10102 8528
rect 9770 8336 9826 8392
rect 9954 8372 9956 8392
rect 9956 8372 10008 8392
rect 10008 8372 10010 8392
rect 9954 8336 10010 8372
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 9770 7948 9826 7984
rect 9770 7928 9772 7948
rect 9772 7928 9824 7948
rect 9824 7928 9826 7948
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 10506 8336 10562 8392
rect 10414 8200 10470 8256
rect 10506 6704 10562 6760
rect 11058 13096 11114 13152
rect 11334 13776 11390 13832
rect 10966 11056 11022 11112
rect 11058 9560 11114 9616
rect 10782 8472 10838 8528
rect 11058 8356 11114 8392
rect 11058 8336 11060 8356
rect 11060 8336 11112 8356
rect 11112 8336 11114 8356
rect 11150 4120 11206 4176
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 11794 12688 11850 12744
rect 11610 8236 11612 8256
rect 11612 8236 11664 8256
rect 11664 8236 11666 8256
rect 11610 8200 11666 8236
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 11886 9152 11942 9208
rect 12254 8880 12310 8936
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 12254 7384 12310 7440
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 12714 11056 12770 11112
rect 12714 9424 12770 9480
rect 13174 12824 13230 12880
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 13266 9152 13322 9208
rect 13174 9036 13230 9072
rect 13174 9016 13176 9036
rect 13176 9016 13228 9036
rect 13228 9016 13230 9036
rect 12990 8916 12992 8936
rect 12992 8916 13044 8936
rect 13044 8916 13046 8936
rect 12990 8880 13046 8916
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 14002 9152 14058 9208
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 14094 7384 14150 7440
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 12898 5364 12954 5400
rect 12898 5344 12900 5364
rect 12900 5344 12952 5364
rect 12952 5344 12954 5364
rect 11978 4800 12034 4856
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 13174 4800 13230 4856
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 14002 5772 14058 5808
rect 14002 5752 14004 5772
rect 14004 5752 14056 5772
rect 14056 5752 14058 5772
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 13542 5072 13598 5128
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 13082 2624 13138 2680
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 15198 9460 15200 9480
rect 15200 9460 15252 9480
rect 15252 9460 15254 9480
rect 15198 9424 15254 9460
rect 15290 9016 15346 9072
rect 16026 5772 16082 5808
rect 16026 5752 16028 5772
rect 16028 5752 16080 5772
rect 16080 5752 16082 5772
rect 15474 5108 15476 5128
rect 15476 5108 15528 5128
rect 15528 5108 15530 5128
rect 15474 5072 15530 5108
rect 16302 6296 16358 6352
rect 16210 5752 16266 5808
rect 16486 6296 16542 6352
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19062 9560 19118 9616
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 13910 856 13966 912
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 10225 18050 10291 18053
rect 10358 18050 10364 18052
rect 10225 18048 10364 18050
rect 10225 17992 10230 18048
rect 10286 17992 10364 18048
rect 10225 17990 10364 17992
rect 10225 17987 10291 17990
rect 10358 17988 10364 17990
rect 10428 17988 10434 18052
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 11329 13834 11395 13837
rect 11462 13834 11468 13836
rect 11329 13832 11468 13834
rect 11329 13776 11334 13832
rect 11390 13776 11468 13832
rect 11329 13774 11468 13776
rect 11329 13771 11395 13774
rect 11462 13772 11468 13774
rect 11532 13772 11538 13836
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 9489 13290 9555 13293
rect 10685 13290 10751 13293
rect 9489 13288 10751 13290
rect 9489 13232 9494 13288
rect 9550 13232 10690 13288
rect 10746 13232 10751 13288
rect 9489 13230 10751 13232
rect 9489 13227 9555 13230
rect 10685 13227 10751 13230
rect 10041 13154 10107 13157
rect 11053 13154 11119 13157
rect 10041 13152 11119 13154
rect 10041 13096 10046 13152
rect 10102 13096 11058 13152
rect 11114 13096 11119 13152
rect 10041 13094 11119 13096
rect 10041 13091 10107 13094
rect 11053 13091 11119 13094
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 10133 13018 10199 13021
rect 10869 13018 10935 13021
rect 10133 13016 10935 13018
rect 10133 12960 10138 13016
rect 10194 12960 10874 13016
rect 10930 12960 10935 13016
rect 10133 12958 10935 12960
rect 10133 12955 10199 12958
rect 10869 12955 10935 12958
rect 9765 12882 9831 12885
rect 13169 12882 13235 12885
rect 9765 12880 13235 12882
rect 9765 12824 9770 12880
rect 9826 12824 13174 12880
rect 13230 12824 13235 12880
rect 9765 12822 13235 12824
rect 9765 12819 9831 12822
rect 13169 12819 13235 12822
rect 9949 12746 10015 12749
rect 10501 12746 10567 12749
rect 9949 12744 10567 12746
rect 9949 12688 9954 12744
rect 10010 12688 10506 12744
rect 10562 12688 10567 12744
rect 9949 12686 10567 12688
rect 9949 12683 10015 12686
rect 10501 12683 10567 12686
rect 11789 12748 11855 12749
rect 11789 12744 11836 12748
rect 11900 12746 11906 12748
rect 11789 12688 11794 12744
rect 11789 12684 11836 12688
rect 11900 12686 11946 12746
rect 11900 12684 11906 12686
rect 11789 12683 11855 12684
rect 10409 12610 10475 12613
rect 10777 12610 10843 12613
rect 10409 12608 10843 12610
rect 10409 12552 10414 12608
rect 10470 12552 10782 12608
rect 10838 12552 10843 12608
rect 10409 12550 10843 12552
rect 10409 12547 10475 12550
rect 10777 12547 10843 12550
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 10358 12276 10364 12340
rect 10428 12338 10434 12340
rect 10777 12338 10843 12341
rect 10428 12336 10843 12338
rect 10428 12280 10782 12336
rect 10838 12280 10843 12336
rect 10428 12278 10843 12280
rect 10428 12276 10434 12278
rect 10777 12275 10843 12278
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 10961 11116 11027 11117
rect 10910 11114 10916 11116
rect 10870 11054 10916 11114
rect 10980 11112 11027 11116
rect 11022 11056 11027 11112
rect 10910 11052 10916 11054
rect 10980 11052 11027 11056
rect 10961 11051 11027 11052
rect 12709 11116 12775 11117
rect 12709 11112 12756 11116
rect 12820 11114 12826 11116
rect 12709 11056 12714 11112
rect 12709 11052 12756 11056
rect 12820 11054 12866 11114
rect 12820 11052 12826 11054
rect 12709 11051 12775 11052
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 5625 10026 5691 10029
rect 8201 10026 8267 10029
rect 5625 10024 8267 10026
rect 5625 9968 5630 10024
rect 5686 9968 8206 10024
rect 8262 9968 8267 10024
rect 5625 9966 8267 9968
rect 5625 9963 5691 9966
rect 8201 9963 8267 9966
rect 4245 9890 4311 9893
rect 6913 9890 6979 9893
rect 4245 9888 6979 9890
rect 4245 9832 4250 9888
rect 4306 9832 6918 9888
rect 6974 9832 6979 9888
rect 4245 9830 6979 9832
rect 4245 9827 4311 9830
rect 6913 9827 6979 9830
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 16896 9759 17212 9760
rect 11053 9618 11119 9621
rect 19057 9618 19123 9621
rect 11053 9616 19123 9618
rect 11053 9560 11058 9616
rect 11114 9560 19062 9616
rect 19118 9560 19123 9616
rect 11053 9558 19123 9560
rect 11053 9555 11119 9558
rect 19057 9555 19123 9558
rect 12709 9482 12775 9485
rect 15193 9482 15259 9485
rect 12709 9480 15259 9482
rect 12709 9424 12714 9480
rect 12770 9424 15198 9480
rect 15254 9424 15259 9480
rect 12709 9422 15259 9424
rect 12709 9419 12775 9422
rect 15193 9419 15259 9422
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 7557 9210 7623 9213
rect 8753 9210 8819 9213
rect 7557 9208 8819 9210
rect 7557 9152 7562 9208
rect 7618 9152 8758 9208
rect 8814 9152 8819 9208
rect 7557 9150 8819 9152
rect 7557 9147 7623 9150
rect 8753 9147 8819 9150
rect 11881 9210 11947 9213
rect 13261 9210 13327 9213
rect 13997 9210 14063 9213
rect 11881 9208 14063 9210
rect 11881 9152 11886 9208
rect 11942 9152 13266 9208
rect 13322 9152 14002 9208
rect 14058 9152 14063 9208
rect 11881 9150 14063 9152
rect 11881 9147 11947 9150
rect 13261 9147 13327 9150
rect 13997 9147 14063 9150
rect 6913 9074 6979 9077
rect 7925 9074 7991 9077
rect 8661 9074 8727 9077
rect 6913 9072 8727 9074
rect 6913 9016 6918 9072
rect 6974 9016 7930 9072
rect 7986 9016 8666 9072
rect 8722 9016 8727 9072
rect 6913 9014 8727 9016
rect 6913 9011 6979 9014
rect 7925 9011 7991 9014
rect 8661 9011 8727 9014
rect 13169 9074 13235 9077
rect 15285 9074 15351 9077
rect 13169 9072 15351 9074
rect 13169 9016 13174 9072
rect 13230 9016 15290 9072
rect 15346 9016 15351 9072
rect 13169 9014 15351 9016
rect 13169 9011 13235 9014
rect 15285 9011 15351 9014
rect 7833 8938 7899 8941
rect 8661 8938 8727 8941
rect 9581 8938 9647 8941
rect 7833 8936 9647 8938
rect 7833 8880 7838 8936
rect 7894 8880 8666 8936
rect 8722 8880 9586 8936
rect 9642 8880 9647 8936
rect 7833 8878 9647 8880
rect 7833 8875 7899 8878
rect 8661 8875 8727 8878
rect 9581 8875 9647 8878
rect 12249 8938 12315 8941
rect 12985 8938 13051 8941
rect 12249 8936 13051 8938
rect 12249 8880 12254 8936
rect 12310 8880 12990 8936
rect 13046 8880 13051 8936
rect 12249 8878 13051 8880
rect 12249 8875 12315 8878
rect 12985 8875 13051 8878
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 10041 8530 10107 8533
rect 10777 8530 10843 8533
rect 10041 8528 10843 8530
rect 10041 8472 10046 8528
rect 10102 8472 10782 8528
rect 10838 8472 10843 8528
rect 10041 8470 10843 8472
rect 10041 8467 10107 8470
rect 10777 8467 10843 8470
rect 9765 8394 9831 8397
rect 9630 8392 9831 8394
rect 9630 8336 9770 8392
rect 9826 8336 9831 8392
rect 9630 8334 9831 8336
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9630 7986 9690 8334
rect 9765 8331 9831 8334
rect 9949 8394 10015 8397
rect 10501 8394 10567 8397
rect 11053 8394 11119 8397
rect 9949 8392 10426 8394
rect 9949 8336 9954 8392
rect 10010 8336 10426 8392
rect 9949 8334 10426 8336
rect 9949 8331 10015 8334
rect 10366 8261 10426 8334
rect 10501 8392 11119 8394
rect 10501 8336 10506 8392
rect 10562 8336 11058 8392
rect 11114 8336 11119 8392
rect 10501 8334 11119 8336
rect 10501 8331 10567 8334
rect 11053 8331 11119 8334
rect 10366 8258 10475 8261
rect 11605 8258 11671 8261
rect 10366 8256 11671 8258
rect 10366 8200 10414 8256
rect 10470 8200 11610 8256
rect 11666 8200 11671 8256
rect 10366 8198 11671 8200
rect 10409 8195 10475 8198
rect 11605 8195 11671 8198
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19253 8127 19569 8128
rect 9765 7986 9831 7989
rect 9630 7984 9831 7986
rect 9630 7928 9770 7984
rect 9826 7928 9831 7984
rect 9630 7926 9831 7928
rect 9765 7923 9831 7926
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 12249 7442 12315 7445
rect 14089 7442 14155 7445
rect 12249 7440 14155 7442
rect 12249 7384 12254 7440
rect 12310 7384 14094 7440
rect 14150 7384 14155 7440
rect 12249 7382 14155 7384
rect 12249 7379 12315 7382
rect 14089 7379 14155 7382
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 7465 6898 7531 6901
rect 8661 6898 8727 6901
rect 7465 6896 8727 6898
rect 7465 6840 7470 6896
rect 7526 6840 8666 6896
rect 8722 6840 8727 6896
rect 7465 6838 8727 6840
rect 7465 6835 7531 6838
rect 8661 6835 8727 6838
rect 4245 6762 4311 6765
rect 10501 6762 10567 6765
rect 4245 6760 10567 6762
rect 4245 6704 4250 6760
rect 4306 6704 10506 6760
rect 10562 6704 10567 6760
rect 4245 6702 10567 6704
rect 4245 6699 4311 6702
rect 10501 6699 10567 6702
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 16297 6354 16363 6357
rect 16481 6354 16547 6357
rect 16297 6352 16547 6354
rect 16297 6296 16302 6352
rect 16358 6296 16486 6352
rect 16542 6296 16547 6352
rect 16297 6294 16547 6296
rect 16297 6291 16363 6294
rect 16481 6291 16547 6294
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 13997 5810 14063 5813
rect 16021 5810 16087 5813
rect 16205 5810 16271 5813
rect 13997 5808 16271 5810
rect 13997 5752 14002 5808
rect 14058 5752 16026 5808
rect 16082 5752 16210 5808
rect 16266 5752 16271 5808
rect 13997 5750 16271 5752
rect 13997 5747 14063 5750
rect 16021 5747 16087 5750
rect 16205 5747 16271 5750
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 12750 5340 12756 5404
rect 12820 5402 12826 5404
rect 12893 5402 12959 5405
rect 12820 5400 12959 5402
rect 12820 5344 12898 5400
rect 12954 5344 12959 5400
rect 12820 5342 12959 5344
rect 12820 5340 12826 5342
rect 12893 5339 12959 5342
rect 6821 5266 6887 5269
rect 8569 5266 8635 5269
rect 6821 5264 8635 5266
rect 6821 5208 6826 5264
rect 6882 5208 8574 5264
rect 8630 5208 8635 5264
rect 6821 5206 8635 5208
rect 6821 5203 6887 5206
rect 8569 5203 8635 5206
rect 13537 5130 13603 5133
rect 15469 5130 15535 5133
rect 13537 5128 15535 5130
rect 13537 5072 13542 5128
rect 13598 5072 15474 5128
rect 15530 5072 15535 5128
rect 13537 5070 15535 5072
rect 13537 5067 13603 5070
rect 15469 5067 15535 5070
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 11973 4858 12039 4861
rect 13169 4858 13235 4861
rect 11973 4856 13235 4858
rect 11973 4800 11978 4856
rect 12034 4800 13174 4856
rect 13230 4800 13235 4856
rect 11973 4798 13235 4800
rect 11973 4795 12039 4798
rect 13169 4795 13235 4798
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 8201 4178 8267 4181
rect 11145 4178 11211 4181
rect 8201 4176 11211 4178
rect 8201 4120 8206 4176
rect 8262 4120 11150 4176
rect 11206 4120 11211 4176
rect 8201 4118 11211 4120
rect 8201 4115 8267 4118
rect 11145 4115 11211 4118
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 11462 2620 11468 2684
rect 11532 2682 11538 2684
rect 13077 2682 13143 2685
rect 11532 2680 13143 2682
rect 11532 2624 13082 2680
rect 13138 2624 13143 2680
rect 11532 2622 13143 2624
rect 11532 2620 11538 2622
rect 13077 2619 13143 2622
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 3877 1458 3943 1461
rect 10910 1458 10916 1460
rect 3877 1456 10916 1458
rect 3877 1400 3882 1456
rect 3938 1400 10916 1456
rect 3877 1398 10916 1400
rect 3877 1395 3943 1398
rect 10910 1396 10916 1398
rect 10980 1396 10986 1460
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 11830 852 11836 916
rect 11900 914 11906 916
rect 13905 914 13971 917
rect 11900 912 13971 914
rect 11900 856 13910 912
rect 13966 856 13971 912
rect 11900 854 13971 856
rect 11900 852 11906 854
rect 13905 851 13971 854
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 10364 17988 10428 18052
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 11468 13772 11532 13836
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 11836 12744 11900 12748
rect 11836 12688 11850 12744
rect 11850 12688 11900 12744
rect 11836 12684 11900 12688
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 10364 12276 10428 12340
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 10916 11112 10980 11116
rect 10916 11056 10966 11112
rect 10966 11056 10980 11112
rect 10916 11052 10980 11056
rect 12756 11112 12820 11116
rect 12756 11056 12770 11112
rect 12770 11056 12820 11112
rect 12756 11052 12820 11056
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 12756 5340 12820 5404
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 11468 2620 11532 2684
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 10916 1396 10980 1460
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 11836 852 11900 916
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 10363 18052 10429 18053
rect 10363 17988 10364 18052
rect 10428 17988 10429 18052
rect 10363 17987 10429 17988
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9821 11456 10141 12480
rect 10366 12341 10426 17987
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 11467 13836 11533 13837
rect 11467 13772 11468 13836
rect 11532 13772 11533 13836
rect 11467 13771 11533 13772
rect 10363 12340 10429 12341
rect 10363 12276 10364 12340
rect 10428 12276 10429 12340
rect 10363 12275 10429 12276
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 10918 1461 10978 11051
rect 11470 2685 11530 13771
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 11835 12748 11901 12749
rect 11835 12684 11836 12748
rect 11900 12684 11901 12748
rect 11835 12683 11901 12684
rect 11467 2684 11533 2685
rect 11467 2620 11468 2684
rect 11532 2620 11533 2684
rect 11467 2619 11533 2620
rect 10915 1460 10981 1461
rect 10915 1396 10916 1460
rect 10980 1396 10981 1460
rect 10915 1395 10981 1396
rect 11838 917 11898 12683
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 12755 11116 12821 11117
rect 12755 11052 12756 11116
rect 12820 11052 12821 11116
rect 12755 11051 12821 11052
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12758 5405 12818 11051
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 12755 5404 12821 5405
rect 12755 5340 12756 5404
rect 12820 5340 12821 5404
rect 12755 5339 12821 5340
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 11835 916 11901 917
rect 11835 852 11836 916
rect 11900 852 11901 916
rect 11835 851 11901 852
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 496 12499 1056
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1720342921
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1720342921
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _286_
timestamp 1720342921
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _287_
timestamp 1720342921
transform 1 0 7636 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_2  _288_
timestamp 1720342921
transform 1 0 9108 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1720342921
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _290_
timestamp 1720342921
transform 1 0 7544 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _291_
timestamp 1720342921
transform 1 0 8372 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _292_
timestamp 1720342921
transform 1 0 7176 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _293_
timestamp 1720342921
transform 1 0 3956 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _294_
timestamp 1720342921
transform 1 0 7360 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _295_
timestamp 1720342921
transform -1 0 10212 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _296_
timestamp 1720342921
transform 1 0 8648 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _297_
timestamp 1720342921
transform 1 0 9200 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _298_
timestamp 1720342921
transform 1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _299_
timestamp 1720342921
transform 1 0 8372 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _300_
timestamp 1720342921
transform 1 0 9016 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _301_
timestamp 1720342921
transform 1 0 9200 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _302_
timestamp 1720342921
transform -1 0 12052 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _303_
timestamp 1720342921
transform 1 0 10304 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _304_
timestamp 1720342921
transform 1 0 9568 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _305_
timestamp 1720342921
transform 1 0 8740 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _306_
timestamp 1720342921
transform 1 0 11684 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _307_
timestamp 1720342921
transform -1 0 11224 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _308_
timestamp 1720342921
transform -1 0 11592 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp 1720342921
transform -1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _310_
timestamp 1720342921
transform -1 0 7636 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _311_
timestamp 1720342921
transform -1 0 9200 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _312_
timestamp 1720342921
transform -1 0 10396 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _313_
timestamp 1720342921
transform -1 0 9660 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _314_
timestamp 1720342921
transform -1 0 8832 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1720342921
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1720342921
transform 1 0 11132 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _317_
timestamp 1720342921
transform -1 0 10488 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _318_
timestamp 1720342921
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _319_
timestamp 1720342921
transform 1 0 9108 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _320_
timestamp 1720342921
transform -1 0 9108 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _321_
timestamp 1720342921
transform -1 0 10120 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _322_
timestamp 1720342921
transform -1 0 9936 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _323_
timestamp 1720342921
transform -1 0 7268 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _324_
timestamp 1720342921
transform 1 0 9844 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _325_
timestamp 1720342921
transform 1 0 14996 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _326_
timestamp 1720342921
transform 1 0 11408 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _327_
timestamp 1720342921
transform 1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _328_
timestamp 1720342921
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _329_
timestamp 1720342921
transform -1 0 11132 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _330_
timestamp 1720342921
transform 1 0 10028 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _331_
timestamp 1720342921
transform -1 0 9384 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _332_
timestamp 1720342921
transform 1 0 6348 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _333_
timestamp 1720342921
transform 1 0 6256 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _334_
timestamp 1720342921
transform -1 0 7084 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _335_
timestamp 1720342921
transform -1 0 9752 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _336_
timestamp 1720342921
transform -1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _337_
timestamp 1720342921
transform 1 0 9476 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _338_
timestamp 1720342921
transform 1 0 7636 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _339_
timestamp 1720342921
transform 1 0 6716 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _340_
timestamp 1720342921
transform -1 0 8832 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _341_
timestamp 1720342921
transform -1 0 7452 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _342_
timestamp 1720342921
transform 1 0 11684 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _343_
timestamp 1720342921
transform -1 0 11316 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _344_
timestamp 1720342921
transform 1 0 11132 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1720342921
transform 1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp 1720342921
transform 1 0 11316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1720342921
transform 1 0 11224 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _348_
timestamp 1720342921
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_2  _349_
timestamp 1720342921
transform 1 0 10948 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp 1720342921
transform -1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _351_
timestamp 1720342921
transform -1 0 7544 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _352_
timestamp 1720342921
transform -1 0 7728 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1720342921
transform -1 0 5612 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _354_
timestamp 1720342921
transform -1 0 11316 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _355_
timestamp 1720342921
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _356_
timestamp 1720342921
transform -1 0 5060 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _357_
timestamp 1720342921
transform 1 0 6072 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _358_
timestamp 1720342921
transform -1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _359_
timestamp 1720342921
transform 1 0 8372 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _360_
timestamp 1720342921
transform -1 0 9292 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _361_
timestamp 1720342921
transform 1 0 7636 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _362_
timestamp 1720342921
transform -1 0 6992 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1720342921
transform -1 0 6992 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1720342921
transform -1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _365_
timestamp 1720342921
transform 1 0 4968 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _366_
timestamp 1720342921
transform 1 0 4692 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _367_
timestamp 1720342921
transform -1 0 4968 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _368_
timestamp 1720342921
transform -1 0 4232 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _369_
timestamp 1720342921
transform -1 0 4692 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _370_
timestamp 1720342921
transform -1 0 5336 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _371_
timestamp 1720342921
transform -1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _372_
timestamp 1720342921
transform 1 0 4600 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _373_
timestamp 1720342921
transform 1 0 3588 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _374_
timestamp 1720342921
transform -1 0 6624 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _375_
timestamp 1720342921
transform -1 0 6900 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _376_
timestamp 1720342921
transform -1 0 7728 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _377_
timestamp 1720342921
transform 1 0 6164 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _378_
timestamp 1720342921
transform 1 0 4048 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _379_
timestamp 1720342921
transform 1 0 3588 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _380_
timestamp 1720342921
transform -1 0 5520 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _381_
timestamp 1720342921
transform 1 0 5796 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _382_
timestamp 1720342921
transform 1 0 4324 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _383_
timestamp 1720342921
transform -1 0 5428 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _384_
timestamp 1720342921
transform -1 0 5612 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1720342921
transform 1 0 3956 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _386_
timestamp 1720342921
transform 1 0 4048 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _387_
timestamp 1720342921
transform 1 0 3404 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _388_
timestamp 1720342921
transform 1 0 7728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _389_
timestamp 1720342921
transform -1 0 6072 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _390_
timestamp 1720342921
transform 1 0 4508 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _391_
timestamp 1720342921
transform 1 0 4876 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _392_
timestamp 1720342921
transform 1 0 6532 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _393_
timestamp 1720342921
transform 1 0 6992 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _394_
timestamp 1720342921
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _395_
timestamp 1720342921
transform -1 0 8096 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _396_
timestamp 1720342921
transform 1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _397_
timestamp 1720342921
transform 1 0 5612 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _398_
timestamp 1720342921
transform 1 0 7268 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _399_
timestamp 1720342921
transform 1 0 7452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _400_
timestamp 1720342921
transform 1 0 8372 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _401_
timestamp 1720342921
transform 1 0 7176 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _402_
timestamp 1720342921
transform -1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _403_
timestamp 1720342921
transform -1 0 8924 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _404_
timestamp 1720342921
transform 1 0 8372 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1720342921
transform -1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _406_
timestamp 1720342921
transform 1 0 10120 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _407_
timestamp 1720342921
transform 1 0 10672 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _408_
timestamp 1720342921
transform 1 0 6808 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _409_
timestamp 1720342921
transform 1 0 7728 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _410_
timestamp 1720342921
transform -1 0 8372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _411_
timestamp 1720342921
transform 1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _412_
timestamp 1720342921
transform 1 0 7452 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _413_
timestamp 1720342921
transform -1 0 7636 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _414_
timestamp 1720342921
transform 1 0 6624 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _415_
timestamp 1720342921
transform 1 0 5888 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1720342921
transform 1 0 6164 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _417_
timestamp 1720342921
transform -1 0 5612 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _418_
timestamp 1720342921
transform -1 0 5612 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _419_
timestamp 1720342921
transform -1 0 5152 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1720342921
transform 1 0 4232 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _421_
timestamp 1720342921
transform -1 0 5428 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _422_
timestamp 1720342921
transform -1 0 5612 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _423_
timestamp 1720342921
transform -1 0 5336 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1720342921
transform 1 0 4324 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _425_
timestamp 1720342921
transform -1 0 5796 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _426_
timestamp 1720342921
transform 1 0 5796 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _427_
timestamp 1720342921
transform -1 0 6440 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1720342921
transform -1 0 4968 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _429_
timestamp 1720342921
transform -1 0 7268 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _430_
timestamp 1720342921
transform 1 0 5888 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _431_
timestamp 1720342921
transform 1 0 6164 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1720342921
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _433_
timestamp 1720342921
transform 1 0 5520 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _434_
timestamp 1720342921
transform 1 0 5704 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _435_
timestamp 1720342921
transform -1 0 5428 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _436_
timestamp 1720342921
transform 1 0 4876 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _437_
timestamp 1720342921
transform 1 0 4232 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1720342921
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _439_
timestamp 1720342921
transform -1 0 3496 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _440_
timestamp 1720342921
transform -1 0 3036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _441_
timestamp 1720342921
transform 1 0 2392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _442_
timestamp 1720342921
transform 1 0 3312 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _443_
timestamp 1720342921
transform 1 0 3220 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _444_
timestamp 1720342921
transform -1 0 4232 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _445_
timestamp 1720342921
transform 1 0 2300 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _446_
timestamp 1720342921
transform -1 0 4416 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _447_
timestamp 1720342921
transform -1 0 3680 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _448_
timestamp 1720342921
transform 1 0 2852 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _449_
timestamp 1720342921
transform -1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1720342921
transform 1 0 13340 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _451_
timestamp 1720342921
transform 1 0 14628 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _452_
timestamp 1720342921
transform 1 0 14168 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 1720342921
transform 1 0 12972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _454_
timestamp 1720342921
transform 1 0 14444 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _455_
timestamp 1720342921
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _456_
timestamp 1720342921
transform -1 0 13524 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 1720342921
transform -1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _458_
timestamp 1720342921
transform 1 0 13524 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _459_
timestamp 1720342921
transform -1 0 12880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _460_
timestamp 1720342921
transform 1 0 12512 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _461_
timestamp 1720342921
transform -1 0 12788 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _462_
timestamp 1720342921
transform 1 0 12144 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _463_
timestamp 1720342921
transform -1 0 17204 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _464_
timestamp 1720342921
transform 1 0 16284 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _465_
timestamp 1720342921
transform 1 0 16560 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _466_
timestamp 1720342921
transform -1 0 15180 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _467_
timestamp 1720342921
transform 1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _468_
timestamp 1720342921
transform -1 0 15364 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _469_
timestamp 1720342921
transform 1 0 11960 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _470_
timestamp 1720342921
transform 1 0 11868 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 1720342921
transform 1 0 11316 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _472_
timestamp 1720342921
transform 1 0 10948 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _473_
timestamp 1720342921
transform -1 0 13800 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _474_
timestamp 1720342921
transform 1 0 15916 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 1720342921
transform -1 0 16008 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1720342921
transform 1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _477_
timestamp 1720342921
transform 1 0 15180 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _478_
timestamp 1720342921
transform 1 0 12880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _479_
timestamp 1720342921
transform 1 0 13708 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _480_
timestamp 1720342921
transform -1 0 13800 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _481_
timestamp 1720342921
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _482_
timestamp 1720342921
transform 1 0 12880 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _483_
timestamp 1720342921
transform 1 0 12880 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _484_
timestamp 1720342921
transform 1 0 13432 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 1720342921
transform 1 0 13800 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _486_
timestamp 1720342921
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _487_
timestamp 1720342921
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _488_
timestamp 1720342921
transform -1 0 17296 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _489_
timestamp 1720342921
transform -1 0 16008 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _490_
timestamp 1720342921
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _491_
timestamp 1720342921
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _492_
timestamp 1720342921
transform 1 0 15180 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _493_
timestamp 1720342921
transform 1 0 16100 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _494_
timestamp 1720342921
transform 1 0 16744 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _495_
timestamp 1720342921
transform 1 0 17020 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _496_
timestamp 1720342921
transform -1 0 17020 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _497_
timestamp 1720342921
transform 1 0 16284 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _498_
timestamp 1720342921
transform -1 0 16836 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _499_
timestamp 1720342921
transform 1 0 14996 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _500_
timestamp 1720342921
transform 1 0 15916 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _501_
timestamp 1720342921
transform -1 0 14904 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _502_
timestamp 1720342921
transform -1 0 14352 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _503_
timestamp 1720342921
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _504_
timestamp 1720342921
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _505_
timestamp 1720342921
transform 1 0 12144 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _506_
timestamp 1720342921
transform 1 0 10120 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _507_
timestamp 1720342921
transform -1 0 16560 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _508_
timestamp 1720342921
transform 1 0 13800 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _509_
timestamp 1720342921
transform -1 0 14260 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _510_
timestamp 1720342921
transform -1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _511_
timestamp 1720342921
transform -1 0 16744 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _512_
timestamp 1720342921
transform 1 0 14260 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _513_
timestamp 1720342921
transform 1 0 15640 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _514_
timestamp 1720342921
transform 1 0 14996 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _515_
timestamp 1720342921
transform -1 0 15180 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _516_
timestamp 1720342921
transform 1 0 14352 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _517_
timestamp 1720342921
transform -1 0 13432 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _518_
timestamp 1720342921
transform 1 0 11592 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _519_
timestamp 1720342921
transform 1 0 10304 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _520_
timestamp 1720342921
transform 1 0 9936 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _521_
timestamp 1720342921
transform -1 0 15824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _522_
timestamp 1720342921
transform -1 0 15640 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _523_
timestamp 1720342921
transform -1 0 14720 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _524_
timestamp 1720342921
transform -1 0 15548 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__o2111ai_1  _525_
timestamp 1720342921
transform 1 0 12604 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1720342921
transform 1 0 12052 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _527_
timestamp 1720342921
transform -1 0 12972 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _528_
timestamp 1720342921
transform 1 0 12144 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _529_
timestamp 1720342921
transform 1 0 10304 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _530_
timestamp 1720342921
transform -1 0 11684 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _531_
timestamp 1720342921
transform 1 0 13524 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _532_
timestamp 1720342921
transform -1 0 14812 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _533_
timestamp 1720342921
transform 1 0 12328 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _534_
timestamp 1720342921
transform 1 0 11684 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _535_
timestamp 1720342921
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _536_
timestamp 1720342921
transform -1 0 11500 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _537_
timestamp 1720342921
transform 1 0 12696 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _538_
timestamp 1720342921
transform 1 0 11960 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _539_
timestamp 1720342921
transform -1 0 12696 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _540_
timestamp 1720342921
transform 1 0 12512 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _541_
timestamp 1720342921
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _542_
timestamp 1720342921
transform -1 0 14168 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _543_
timestamp 1720342921
transform -1 0 16744 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _544_
timestamp 1720342921
transform 1 0 13984 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _545_
timestamp 1720342921
transform -1 0 13984 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _546_
timestamp 1720342921
transform 1 0 12972 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _547_
timestamp 1720342921
transform -1 0 14628 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _548_
timestamp 1720342921
transform -1 0 14168 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _549_
timestamp 1720342921
transform -1 0 13984 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _550_
timestamp 1720342921
transform 1 0 10948 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _551_
timestamp 1720342921
transform 1 0 11316 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _552_
timestamp 1720342921
transform 1 0 11684 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _553_
timestamp 1720342921
transform -1 0 13248 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _554_
timestamp 1720342921
transform 1 0 10212 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _555_
timestamp 1720342921
transform 1 0 9936 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _556_
timestamp 1720342921
transform -1 0 8004 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _557_
timestamp 1720342921
transform 1 0 9936 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _558_
timestamp 1720342921
transform 1 0 8096 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _559_
timestamp 1720342921
transform -1 0 8556 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _560_
timestamp 1720342921
transform 1 0 8372 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _561_
timestamp 1720342921
transform 1 0 6256 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _562_
timestamp 1720342921
transform 1 0 5796 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _563_
timestamp 1720342921
transform 1 0 3680 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _564_
timestamp 1720342921
transform 1 0 3680 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _565_
timestamp 1720342921
transform 1 0 4968 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _566_
timestamp 1720342921
transform 1 0 6808 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _567_
timestamp 1720342921
transform 1 0 5796 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _568_
timestamp 1720342921
transform 1 0 3772 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _569_
timestamp 1720342921
transform 1 0 2208 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _570_
timestamp 1720342921
transform 1 0 1840 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _571_
timestamp 1720342921
transform 1 0 2300 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _572_
timestamp 1720342921
transform -1 0 4048 0 -1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _573_
timestamp 1720342921
transform -1 0 14260 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _574_
timestamp 1720342921
transform -1 0 13248 0 -1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _575_
timestamp 1720342921
transform -1 0 9200 0 -1 2720
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _576_
timestamp 1720342921
transform 1 0 10028 0 1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _577_
timestamp 1720342921
transform 1 0 13248 0 -1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _578_
timestamp 1720342921
transform 1 0 13616 0 1 544
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _579_
timestamp 1720342921
transform 1 0 16468 0 -1 1632
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _580__12
timestamp 1720342921
transform 1 0 15180 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _580_
timestamp 1720342921
transform 1 0 14812 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_2  _581_
timestamp 1720342921
transform 1 0 8464 0 -1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _582_
timestamp 1720342921
transform 1 0 9384 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _583_
timestamp 1720342921
transform 1 0 8556 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _584_
timestamp 1720342921
transform 1 0 2852 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _585_
timestamp 1720342921
transform 1 0 8464 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _586_
timestamp 1720342921
transform 1 0 9292 0 1 3808
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _587_
timestamp 1720342921
transform 1 0 14352 0 1 11424
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _588_
timestamp 1720342921
transform 1 0 13616 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _589_
timestamp 1720342921
transform 1 0 11960 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _590_
timestamp 1720342921
transform 1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _591_
timestamp 1720342921
transform -1 0 13340 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _592_
timestamp 1720342921
transform -1 0 11868 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _593_
timestamp 1720342921
transform -1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _594_
timestamp 1720342921
transform 1 0 6716 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _595_
timestamp 1720342921
transform -1 0 12420 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _596_
timestamp 1720342921
transform 1 0 8648 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _597_
timestamp 1720342921
transform 1 0 10212 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _598_
timestamp 1720342921
transform 1 0 6808 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _599_
timestamp 1720342921
transform 1 0 3864 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _600_
timestamp 1720342921
transform -1 0 3772 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _601_
timestamp 1720342921
transform 1 0 5796 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _602_
timestamp 1720342921
transform 1 0 10856 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _603_
timestamp 1720342921
transform 1 0 10948 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1720342921
transform -1 0 2300 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1720342921
transform -1 0 11132 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1720342921
transform 1 0 8372 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1720342921
transform 1 0 10948 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1720342921
transform -1 0 9108 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1720342921
transform 1 0 10948 0 -1 13600
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1720342921
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1720342921
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1720342921
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1720342921
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1720342921
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 1720342921
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1720342921
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1720342921
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1720342921
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1720342921
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1720342921
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1720342921
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1720342921
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1720342921
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1720342921
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1720342921
transform 1 0 13524 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_159
timestamp 1720342921
transform 1 0 15180 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1720342921
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1720342921
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1720342921
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1720342921
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197
timestamp 1720342921
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_201
timestamp 1720342921
transform 1 0 19044 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1720342921
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_15
timestamp 1720342921
transform 1 0 1932 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_19
timestamp 1720342921
transform 1 0 2300 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_38
timestamp 1720342921
transform 1 0 4048 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_50
timestamp 1720342921
transform 1 0 5152 0 -1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1720342921
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1720342921
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1720342921
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1720342921
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1720342921
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1720342921
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1720342921
transform 1 0 10948 0 -1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_155
timestamp 1720342921
transform 1 0 14812 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1720342921
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_169
timestamp 1720342921
transform 1 0 16100 0 -1 1632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_190
timestamp 1720342921
transform 1 0 18032 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1720342921
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1720342921
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1720342921
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1720342921
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1720342921
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1720342921
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1720342921
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1720342921
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1720342921
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1720342921
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_97
timestamp 1720342921
transform 1 0 9476 0 1 1632
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_120
timestamp 1720342921
transform 1 0 11592 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_132
timestamp 1720342921
transform 1 0 12696 0 1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1720342921
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1720342921
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1720342921
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1720342921
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1720342921
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1720342921
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1720342921
transform 1 0 18676 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1720342921
transform 1 0 19044 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1720342921
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1720342921
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1720342921
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1720342921
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1720342921
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1720342921
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1720342921
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1720342921
transform 1 0 6900 0 -1 2720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_94
timestamp 1720342921
transform 1 0 9200 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_106
timestamp 1720342921
transform 1 0 10304 0 -1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1720342921
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_125
timestamp 1720342921
transform 1 0 12052 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_131
timestamp 1720342921
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1720342921
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1720342921
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1720342921
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1720342921
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1720342921
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_193
timestamp 1720342921
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 1720342921
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1720342921
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1720342921
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1720342921
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1720342921
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1720342921
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1720342921
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1720342921
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1720342921
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1720342921
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1720342921
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1720342921
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1720342921
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1720342921
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1720342921
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1720342921
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1720342921
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1720342921
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1720342921
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1720342921
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1720342921
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1720342921
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1720342921
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1720342921
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1720342921
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1720342921
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1720342921
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1720342921
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1720342921
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1720342921
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1720342921
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1720342921
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_81
timestamp 1720342921
transform 1 0 8004 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_85
timestamp 1720342921
transform 1 0 8372 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1720342921
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1720342921
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_129
timestamp 1720342921
transform 1 0 12420 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_141
timestamp 1720342921
transform 1 0 13524 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_153
timestamp 1720342921
transform 1 0 14628 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1720342921
transform 1 0 15732 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1720342921
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1720342921
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1720342921
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1720342921
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1720342921
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1720342921
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1720342921
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1720342921
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1720342921
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_53
timestamp 1720342921
transform 1 0 5428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 1720342921
transform 1 0 7268 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1720342921
transform 1 0 8004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_91
timestamp 1720342921
transform 1 0 8924 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1720342921
transform 1 0 13064 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_148
timestamp 1720342921
transform 1 0 14168 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_154
timestamp 1720342921
transform 1 0 14720 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_166
timestamp 1720342921
transform 1 0 15824 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_178
timestamp 1720342921
transform 1 0 16928 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_190
timestamp 1720342921
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1720342921
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1720342921
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1720342921
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1720342921
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1720342921
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1720342921
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1720342921
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1720342921
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_57
timestamp 1720342921
transform 1 0 5796 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_63
timestamp 1720342921
transform 1 0 6348 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_71
timestamp 1720342921
transform 1 0 7084 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_91
timestamp 1720342921
transform 1 0 8924 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1720342921
transform 1 0 10028 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1720342921
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1720342921
transform 1 0 11316 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_130
timestamp 1720342921
transform 1 0 12512 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_138
timestamp 1720342921
transform 1 0 13248 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1720342921
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1720342921
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1720342921
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp 1720342921
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_201
timestamp 1720342921
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1720342921
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1720342921
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1720342921
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1720342921
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1720342921
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_53
timestamp 1720342921
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_63
timestamp 1720342921
transform 1 0 6348 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_92
timestamp 1720342921
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_104
timestamp 1720342921
transform 1 0 10120 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_112
timestamp 1720342921
transform 1 0 10856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_120
timestamp 1720342921
transform 1 0 11592 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1720342921
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1720342921
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1720342921
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_164
timestamp 1720342921
transform 1 0 15640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_168
timestamp 1720342921
transform 1 0 16008 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_174
timestamp 1720342921
transform 1 0 16560 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_186
timestamp 1720342921
transform 1 0 17664 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1720342921
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_197
timestamp 1720342921
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_201
timestamp 1720342921
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1720342921
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_15
timestamp 1720342921
transform 1 0 1932 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_23
timestamp 1720342921
transform 1 0 2668 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_41
timestamp 1720342921
transform 1 0 4324 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_77
timestamp 1720342921
transform 1 0 7636 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_89
timestamp 1720342921
transform 1 0 8740 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_140
timestamp 1720342921
transform 1 0 13432 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_147
timestamp 1720342921
transform 1 0 14076 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_151
timestamp 1720342921
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_155
timestamp 1720342921
transform 1 0 14812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1720342921
transform 1 0 15180 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1720342921
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_179
timestamp 1720342921
transform 1 0 17020 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_191
timestamp 1720342921
transform 1 0 18124 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_199
timestamp 1720342921
transform 1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1720342921
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1720342921
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1720342921
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1720342921
transform 1 0 3220 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_46
timestamp 1720342921
transform 1 0 4784 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_60
timestamp 1720342921
transform 1 0 6072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_72
timestamp 1720342921
transform 1 0 7176 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_124
timestamp 1720342921
transform 1 0 11960 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_136
timestamp 1720342921
transform 1 0 13064 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_149
timestamp 1720342921
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_157
timestamp 1720342921
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_184
timestamp 1720342921
transform 1 0 17480 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1720342921
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1720342921
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1720342921
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1720342921
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1720342921
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_39
timestamp 1720342921
transform 1 0 4140 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1720342921
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1720342921
transform 1 0 6900 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_78
timestamp 1720342921
transform 1 0 7728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_103
timestamp 1720342921
transform 1 0 10028 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_107
timestamp 1720342921
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_116
timestamp 1720342921
transform 1 0 11224 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_122
timestamp 1720342921
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_127
timestamp 1720342921
transform 1 0 12236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_134
timestamp 1720342921
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_141
timestamp 1720342921
transform 1 0 13524 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_153
timestamp 1720342921
transform 1 0 14628 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1720342921
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1720342921
transform 1 0 15916 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_174
timestamp 1720342921
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_186
timestamp 1720342921
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_198
timestamp 1720342921
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1720342921
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1720342921
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1720342921
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1720342921
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_38
timestamp 1720342921
transform 1 0 4048 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_44
timestamp 1720342921
transform 1 0 4600 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_50
timestamp 1720342921
transform 1 0 5152 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_54
timestamp 1720342921
transform 1 0 5520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_58
timestamp 1720342921
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_62
timestamp 1720342921
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_66
timestamp 1720342921
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_71
timestamp 1720342921
transform 1 0 7084 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1720342921
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_88
timestamp 1720342921
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1720342921
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_112
timestamp 1720342921
transform 1 0 10856 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_119
timestamp 1720342921
transform 1 0 11500 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1720342921
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_145
timestamp 1720342921
transform 1 0 13892 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_156
timestamp 1720342921
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_162
timestamp 1720342921
transform 1 0 15456 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_170
timestamp 1720342921
transform 1 0 16192 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1720342921
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1720342921
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1720342921
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1720342921
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1720342921
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1720342921
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1720342921
transform 1 0 1932 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_35
timestamp 1720342921
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_40
timestamp 1720342921
transform 1 0 4232 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1720342921
transform 1 0 5520 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_70
timestamp 1720342921
transform 1 0 6992 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_82
timestamp 1720342921
transform 1 0 8096 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_94
timestamp 1720342921
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 1720342921
transform 1 0 10396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1720342921
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1720342921
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 1720342921
transform 1 0 12052 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 1720342921
transform 1 0 12420 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_141
timestamp 1720342921
transform 1 0 13524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_153
timestamp 1720342921
transform 1 0 14628 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_163
timestamp 1720342921
transform 1 0 15548 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_182
timestamp 1720342921
transform 1 0 17296 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_194
timestamp 1720342921
transform 1 0 18400 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1720342921
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1720342921
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1720342921
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1720342921
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_55
timestamp 1720342921
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_66
timestamp 1720342921
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1720342921
transform 1 0 7268 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1720342921
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1720342921
transform 1 0 8372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_104
timestamp 1720342921
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_125
timestamp 1720342921
transform 1 0 12052 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1720342921
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_149
timestamp 1720342921
transform 1 0 14260 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_156
timestamp 1720342921
transform 1 0 14904 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_162
timestamp 1720342921
transform 1 0 15456 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_166
timestamp 1720342921
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_176
timestamp 1720342921
transform 1 0 16744 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1720342921
transform 1 0 17848 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1720342921
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1720342921
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1720342921
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1720342921
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1720342921
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1720342921
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1720342921
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1720342921
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1720342921
transform 1 0 5796 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp 1720342921
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_95
timestamp 1720342921
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_103
timestamp 1720342921
transform 1 0 10028 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1720342921
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1720342921
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_123
timestamp 1720342921
transform 1 0 11868 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_129
timestamp 1720342921
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_133
timestamp 1720342921
transform 1 0 12788 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_150
timestamp 1720342921
transform 1 0 14352 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_158
timestamp 1720342921
transform 1 0 15088 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_164
timestamp 1720342921
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1720342921
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1720342921
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_193
timestamp 1720342921
transform 1 0 18308 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_201
timestamp 1720342921
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1720342921
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1720342921
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1720342921
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1720342921
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_41
timestamp 1720342921
transform 1 0 4324 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_51
timestamp 1720342921
transform 1 0 5244 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_59
timestamp 1720342921
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_69
timestamp 1720342921
transform 1 0 6900 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_78
timestamp 1720342921
transform 1 0 7728 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1720342921
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_122
timestamp 1720342921
transform 1 0 11776 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1720342921
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_149
timestamp 1720342921
transform 1 0 14260 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_178
timestamp 1720342921
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_190
timestamp 1720342921
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1720342921
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1720342921
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1720342921
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1720342921
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_27
timestamp 1720342921
transform 1 0 3036 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1720342921
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1720342921
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_61
timestamp 1720342921
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_68
timestamp 1720342921
transform 1 0 6808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_76
timestamp 1720342921
transform 1 0 7544 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_84
timestamp 1720342921
transform 1 0 8280 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_90
timestamp 1720342921
transform 1 0 8832 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_94
timestamp 1720342921
transform 1 0 9200 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_106
timestamp 1720342921
transform 1 0 10304 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_121
timestamp 1720342921
transform 1 0 11684 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_132
timestamp 1720342921
transform 1 0 12696 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_147
timestamp 1720342921
transform 1 0 14076 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1720342921
transform 1 0 15640 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_172
timestamp 1720342921
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_184
timestamp 1720342921
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_196
timestamp 1720342921
transform 1 0 18584 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1720342921
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1720342921
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1720342921
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1720342921
transform 1 0 3220 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1720342921
transform 1 0 3956 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_45
timestamp 1720342921
transform 1 0 4692 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_55
timestamp 1720342921
transform 1 0 5612 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_61
timestamp 1720342921
transform 1 0 6164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1720342921
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_85
timestamp 1720342921
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_99
timestamp 1720342921
transform 1 0 9660 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_118
timestamp 1720342921
transform 1 0 11408 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1720342921
transform 1 0 12512 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1720342921
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1720342921
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_153
timestamp 1720342921
transform 1 0 14628 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_171
timestamp 1720342921
transform 1 0 16284 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_183
timestamp 1720342921
transform 1 0 17388 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1720342921
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1720342921
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1720342921
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1720342921
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1720342921
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 1720342921
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_35
timestamp 1720342921
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1720342921
transform 1 0 5336 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1720342921
transform 1 0 5796 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1720342921
transform 1 0 6900 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_81
timestamp 1720342921
transform 1 0 8004 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_85
timestamp 1720342921
transform 1 0 8372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1720342921
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1720342921
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_129
timestamp 1720342921
transform 1 0 12420 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_137
timestamp 1720342921
transform 1 0 13156 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_147
timestamp 1720342921
transform 1 0 14076 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_153
timestamp 1720342921
transform 1 0 14628 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1720342921
transform 1 0 15732 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1720342921
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1720342921
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_193
timestamp 1720342921
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp 1720342921
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1720342921
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1720342921
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1720342921
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1720342921
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1720342921
transform 1 0 4324 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 1720342921
transform 1 0 5428 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_62
timestamp 1720342921
transform 1 0 6256 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1720342921
transform 1 0 8372 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_93
timestamp 1720342921
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_100
timestamp 1720342921
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_112
timestamp 1720342921
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_129
timestamp 1720342921
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_149
timestamp 1720342921
transform 1 0 14260 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_167
timestamp 1720342921
transform 1 0 15916 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_179
timestamp 1720342921
transform 1 0 17020 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_191
timestamp 1720342921
transform 1 0 18124 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1720342921
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1720342921
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1720342921
transform 1 0 19044 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1720342921
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_15
timestamp 1720342921
transform 1 0 1932 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_34
timestamp 1720342921
transform 1 0 3680 0 -1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_43
timestamp 1720342921
transform 1 0 4508 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1720342921
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_76
timestamp 1720342921
transform 1 0 7544 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_88
timestamp 1720342921
transform 1 0 8648 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_100
timestamp 1720342921
transform 1 0 9752 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1720342921
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_153
timestamp 1720342921
transform 1 0 14628 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1720342921
transform 1 0 15732 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1720342921
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1720342921
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 1720342921
transform 1 0 18308 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1720342921
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1720342921
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1720342921
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1720342921
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_29
timestamp 1720342921
transform 1 0 3220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_51
timestamp 1720342921
transform 1 0 5244 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1720342921
transform 1 0 8372 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_97
timestamp 1720342921
transform 1 0 9476 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_113
timestamp 1720342921
transform 1 0 10948 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_121
timestamp 1720342921
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_130
timestamp 1720342921
transform 1 0 12512 0 1 12512
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1720342921
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1720342921
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1720342921
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1720342921
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1720342921
transform 1 0 17940 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1720342921
transform 1 0 18492 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1720342921
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1720342921
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1720342921
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_15
timestamp 1720342921
transform 1 0 1932 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_19
timestamp 1720342921
transform 1 0 2300 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1720342921
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1720342921
transform 1 0 5796 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_93
timestamp 1720342921
transform 1 0 9108 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_102
timestamp 1720342921
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1720342921
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_133
timestamp 1720342921
transform 1 0 12788 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_139
timestamp 1720342921
transform 1 0 13340 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_148
timestamp 1720342921
transform 1 0 14168 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1720342921
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1720342921
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1720342921
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_193
timestamp 1720342921
transform 1 0 18308 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1720342921
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1720342921
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_15
timestamp 1720342921
transform 1 0 1932 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_22
timestamp 1720342921
transform 1 0 2576 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_32
timestamp 1720342921
transform 1 0 3496 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_36
timestamp 1720342921
transform 1 0 3864 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_43
timestamp 1720342921
transform 1 0 4508 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_47
timestamp 1720342921
transform 1 0 4876 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_53
timestamp 1720342921
transform 1 0 5428 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_57
timestamp 1720342921
transform 1 0 5796 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_63
timestamp 1720342921
transform 1 0 6348 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_71
timestamp 1720342921
transform 1 0 7084 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_75
timestamp 1720342921
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_104
timestamp 1720342921
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1720342921
transform 1 0 11224 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1720342921
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_158
timestamp 1720342921
transform 1 0 15088 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_170
timestamp 1720342921
transform 1 0 16192 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_182
timestamp 1720342921
transform 1 0 17296 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1720342921
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1720342921
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_201
timestamp 1720342921
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_3
timestamp 1720342921
transform 1 0 828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_11
timestamp 1720342921
transform 1 0 1564 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_40
timestamp 1720342921
transform 1 0 4232 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_52
timestamp 1720342921
transform 1 0 5336 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_64
timestamp 1720342921
transform 1 0 6440 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_72
timestamp 1720342921
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_97
timestamp 1720342921
transform 1 0 9476 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_101
timestamp 1720342921
transform 1 0 9844 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1720342921
transform 1 0 10212 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1720342921
transform 1 0 10764 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_121
timestamp 1720342921
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_133
timestamp 1720342921
transform 1 0 12788 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1720342921
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1720342921
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1720342921
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_193
timestamp 1720342921
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_201
timestamp 1720342921
transform 1 0 19044 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1720342921
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_15
timestamp 1720342921
transform 1 0 1932 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_23
timestamp 1720342921
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_34
timestamp 1720342921
transform 1 0 3680 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_42
timestamp 1720342921
transform 1 0 4416 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_64
timestamp 1720342921
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1720342921
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_90
timestamp 1720342921
transform 1 0 8832 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_102
timestamp 1720342921
transform 1 0 9936 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_114
timestamp 1720342921
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_119
timestamp 1720342921
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_125
timestamp 1720342921
transform 1 0 12052 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1720342921
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1720342921
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_146
timestamp 1720342921
transform 1 0 13984 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_158
timestamp 1720342921
transform 1 0 15088 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_170
timestamp 1720342921
transform 1 0 16192 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_182
timestamp 1720342921
transform 1 0 17296 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1720342921
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1720342921
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp 1720342921
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1720342921
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_15
timestamp 1720342921
transform 1 0 1932 0 -1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_42
timestamp 1720342921
transform 1 0 4416 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1720342921
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_62
timestamp 1720342921
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_89
timestamp 1720342921
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_100
timestamp 1720342921
transform 1 0 9752 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1720342921
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1720342921
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1720342921
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1720342921
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1720342921
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1720342921
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1720342921
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_193
timestamp 1720342921
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_201
timestamp 1720342921
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1720342921
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1720342921
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1720342921
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1720342921
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_44
timestamp 1720342921
transform 1 0 4600 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_57
timestamp 1720342921
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_65
timestamp 1720342921
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1720342921
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_92
timestamp 1720342921
transform 1 0 9016 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_105
timestamp 1720342921
transform 1 0 10212 0 1 15776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_144
timestamp 1720342921
transform 1 0 13800 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_156
timestamp 1720342921
transform 1 0 14904 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_168
timestamp 1720342921
transform 1 0 16008 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_180
timestamp 1720342921
transform 1 0 17112 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1720342921
transform 1 0 18216 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1720342921
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1720342921
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1720342921
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1720342921
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_27
timestamp 1720342921
transform 1 0 3036 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_33
timestamp 1720342921
transform 1 0 3588 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1720342921
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1720342921
transform 1 0 5796 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_61
timestamp 1720342921
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_92
timestamp 1720342921
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1720342921
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_145
timestamp 1720342921
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_157
timestamp 1720342921
transform 1 0 14996 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1720342921
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1720342921
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1720342921
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp 1720342921
transform 1 0 18308 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1720342921
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1720342921
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1720342921
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1720342921
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1720342921
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_41
timestamp 1720342921
transform 1 0 4324 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_47
timestamp 1720342921
transform 1 0 4876 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1720342921
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1720342921
transform 1 0 6532 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_77
timestamp 1720342921
transform 1 0 7636 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1720342921
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_91
timestamp 1720342921
transform 1 0 8924 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_103
timestamp 1720342921
transform 1 0 10028 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_117
timestamp 1720342921
transform 1 0 11316 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1720342921
transform 1 0 13064 0 1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1720342921
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_153
timestamp 1720342921
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_176
timestamp 1720342921
transform 1 0 16744 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_188
timestamp 1720342921
transform 1 0 17848 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1720342921
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1720342921
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1720342921
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1720342921
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1720342921
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_39
timestamp 1720342921
transform 1 0 4140 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1720342921
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1720342921
transform 1 0 5796 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_65
timestamp 1720342921
transform 1 0 6532 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_77
timestamp 1720342921
transform 1 0 7636 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_81
timestamp 1720342921
transform 1 0 8004 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_85
timestamp 1720342921
transform 1 0 8372 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_95
timestamp 1720342921
transform 1 0 9292 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_103
timestamp 1720342921
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_121
timestamp 1720342921
transform 1 0 11684 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_138
timestamp 1720342921
transform 1 0 13248 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_150
timestamp 1720342921
transform 1 0 14352 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_158
timestamp 1720342921
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 1720342921
transform 1 0 15456 0 -1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1720342921
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1720342921
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1720342921
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_201
timestamp 1720342921
transform 1 0 19044 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1720342921
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1720342921
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1720342921
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_29
timestamp 1720342921
transform 1 0 3220 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_33
timestamp 1720342921
transform 1 0 3588 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_55
timestamp 1720342921
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_73
timestamp 1720342921
transform 1 0 7268 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_101
timestamp 1720342921
transform 1 0 9844 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1720342921
transform 1 0 13340 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1720342921
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1720342921
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_165
timestamp 1720342921
transform 1 0 15732 0 1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_176
timestamp 1720342921
transform 1 0 16744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_188
timestamp 1720342921
transform 1 0 17848 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1720342921
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1720342921
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1720342921
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_8
timestamp 1720342921
transform 1 0 1288 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_20
timestamp 1720342921
transform 1 0 2392 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp 1720342921
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_29
timestamp 1720342921
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_37
timestamp 1720342921
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp 1720342921
transform 1 0 4508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1720342921
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1720342921
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_64
timestamp 1720342921
transform 1 0 6440 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_79
timestamp 1720342921
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp 1720342921
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_85
timestamp 1720342921
transform 1 0 8372 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_93
timestamp 1720342921
transform 1 0 9108 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1720342921
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1720342921
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_116
timestamp 1720342921
transform 1 0 11224 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_124
timestamp 1720342921
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_129
timestamp 1720342921
transform 1 0 12420 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_133
timestamp 1720342921
transform 1 0 12788 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1720342921
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_141
timestamp 1720342921
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_147
timestamp 1720342921
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1720342921
transform 1 0 14444 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1720342921
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1720342921
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_172
timestamp 1720342921
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_187
timestamp 1720342921
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1720342921
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1720342921
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1720342921
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1720342921
transform -1 0 9476 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1720342921
transform -1 0 11684 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1720342921
transform -1 0 8740 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1720342921
transform -1 0 11316 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1720342921
transform -1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1720342921
transform 1 0 11868 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1720342921
transform -1 0 13064 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1720342921
transform -1 0 13156 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1720342921
transform -1 0 4232 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1720342921
transform -1 0 8464 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1720342921
transform -1 0 7452 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1720342921
transform -1 0 15824 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1720342921
transform -1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1720342921
transform -1 0 16376 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1720342921
transform -1 0 14444 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1720342921
transform -1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1720342921
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1720342921
transform 1 0 9200 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1720342921
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1720342921
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1720342921
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1720342921
transform 1 0 2576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1720342921
transform 1 0 920 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1720342921
transform 1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1720342921
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1720342921
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1720342921
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1720342921
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1720342921
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1720342921
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1720342921
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1720342921
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1720342921
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1720342921
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1720342921
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1720342921
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1720342921
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1720342921
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1720342921
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1720342921
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1720342921
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1720342921
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1720342921
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1720342921
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1720342921
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1720342921
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1720342921
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1720342921
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1720342921
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1720342921
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1720342921
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1720342921
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1720342921
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1720342921
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1720342921
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1720342921
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1720342921
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1720342921
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1720342921
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1720342921
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1720342921
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1720342921
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1720342921
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1720342921
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1720342921
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1720342921
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1720342921
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1720342921
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1720342921
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1720342921
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1720342921
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1720342921
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1720342921
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1720342921
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1720342921
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1720342921
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1720342921
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1720342921
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1720342921
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1720342921
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1720342921
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1720342921
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1720342921
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1720342921
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1720342921
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1720342921
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1720342921
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1720342921
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1720342921
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1720342921
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1720342921
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1720342921
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp 1720342921
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1720342921
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1720342921
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1720342921
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1720342921
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1720342921
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1720342921
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1720342921
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1720342921
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1720342921
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1720342921
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1720342921
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1720342921
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1720342921
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1720342921
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1720342921
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1720342921
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1720342921
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1720342921
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1720342921
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1720342921
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1720342921
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1720342921
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1720342921
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1720342921
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1720342921
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1720342921
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1720342921
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1720342921
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1720342921
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1720342921
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1720342921
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1720342921
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1720342921
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1720342921
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1720342921
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1720342921
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1720342921
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1720342921
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1720342921
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1720342921
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1720342921
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1720342921
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1720342921
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1720342921
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1720342921
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1720342921
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1720342921
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1720342921
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1720342921
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1720342921
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1720342921
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1720342921
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1720342921
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1720342921
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1720342921
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1720342921
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1720342921
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1720342921
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1720342921
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1720342921
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1720342921
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1720342921
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1720342921
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1720342921
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1720342921
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1720342921
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1720342921
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1720342921
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1720342921
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1720342921
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1720342921
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1720342921
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1720342921
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1720342921
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1720342921
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1720342921
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1720342921
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1720342921
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1720342921
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1720342921
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1720342921
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1720342921
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1720342921
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1720342921
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1720342921
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1720342921
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1720342921
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1720342921
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1720342921
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1720342921
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1720342921
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1720342921
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1720342921
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1720342921
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1720342921
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1720342921
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1720342921
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1720342921
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1720342921
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1720342921
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1720342921
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1720342921
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1720342921
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1720342921
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1720342921
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1720342921
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1720342921
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1720342921
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1720342921
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1720342921
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1720342921
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1720342921
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1720342921
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1720342921
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1720342921
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1720342921
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1720342921
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1720342921
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1720342921
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1720342921
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1720342921
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1720342921
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1720342921
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1720342921
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1720342921
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 10061 19040 10061 19040 4 VGND
rlabel metal1 s 9982 18496 9982 18496 4 VPWR
rlabel metal2 s 6946 11186 6946 11186 4 _000_
rlabel metal1 s 4048 10778 4048 10778 4 _001_
rlabel metal2 s 3450 7718 3450 7718 4 _002_
rlabel metal1 s 5872 3978 5872 3978 4 _003_
rlabel metal2 s 8234 4301 8234 4301 4 _004_
rlabel metal1 s 11168 3570 11168 3570 4 _005_
rlabel metal1 s 12374 11220 12374 11220 4 _006_
rlabel metal2 s 13846 11662 13846 11662 4 _007_
rlabel metal2 s 14030 8024 14030 8024 4 _008_
rlabel metal2 s 13018 4556 13018 4556 4 _009_
rlabel metal1 s 12144 4250 12144 4250 4 _010_
rlabel metal2 s 12834 3876 12834 3876 4 _011_
rlabel metal2 s 11638 6630 11638 6630 4 _012_
rlabel metal1 s 16429 17102 16429 17102 4 _013_
rlabel metal1 s 8418 17850 8418 17850 4 _014_
rlabel metal1 s 7452 16014 7452 16014 4 _015_
rlabel metal2 s 6113 18122 6113 18122 4 _016_
rlabel metal2 s 4278 17986 4278 17986 4 _017_
rlabel metal2 s 4370 16422 4370 16422 4 _018_
rlabel metal1 s 5090 14858 5090 14858 4 _019_
rlabel metal1 s 7217 12682 7217 12682 4 _020_
rlabel metal2 s 5750 12070 5750 12070 4 _021_
rlabel metal1 s 4181 12682 4181 12682 4 _022_
rlabel metal2 s 2525 12274 2525 12274 4 _023_
rlabel metal1 s 2254 14042 2254 14042 4 _024_
rlabel metal1 s 3128 15130 3128 15130 4 _025_
rlabel metal1 s 3828 1394 3828 1394 4 _026_
rlabel metal1 s 14551 2550 14551 2550 4 _027_
rlabel metal1 s 12332 1462 12332 1462 4 _028_
rlabel metal1 s 9583 2550 9583 2550 4 _029_
rlabel metal1 s 10483 1802 10483 1802 4 _030_
rlabel metal3 s 12305 2652 12305 2652 4 _031_
rlabel metal3 s 12903 884 12903 884 4 _032_
rlabel metal1 s 16744 1530 16744 1530 4 _033_
rlabel metal1 s 5796 7310 5796 7310 4 _034_
rlabel metal1 s 6210 8806 6210 8806 4 _035_
rlabel metal1 s 8234 5168 8234 5168 4 _036_
rlabel metal1 s 7222 4624 7222 4624 4 _037_
rlabel metal1 s 8556 5134 8556 5134 4 _038_
rlabel metal1 s 8924 5134 8924 5134 4 _039_
rlabel metal1 s 14536 11322 14536 11322 4 _040_
rlabel metal2 s 13933 14450 13933 14450 4 _041_
rlabel metal1 s 12082 15946 12082 15946 4 _042_
rlabel metal2 s 12374 17000 12374 17000 4 _043_
rlabel metal2 s 12650 17986 12650 17986 4 _044_
rlabel metal1 s 10948 17850 10948 17850 4 _045_
rlabel metal1 s 11412 16694 11412 16694 4 _046_
rlabel metal1 s 7217 14926 7217 14926 4 _047_
rlabel metal1 s 11320 15606 11320 15606 4 _048_
rlabel metal2 s 8965 13770 8965 13770 4 _049_
rlabel metal1 s 10432 6222 10432 6222 4 _050_
rlabel metal2 s 7314 14212 7314 14212 4 _051_
rlabel metal2 s 4462 14212 4462 14212 4 _052_
rlabel metal2 s 9246 13804 9246 13804 4 _053_
rlabel metal1 s 9982 16218 9982 16218 4 _054_
rlabel metal2 s 9246 17068 9246 17068 4 _055_
rlabel metal1 s 9614 13294 9614 13294 4 _056_
rlabel metal1 s 9062 16558 9062 16558 4 _057_
rlabel metal2 s 9062 15810 9062 15810 4 _058_
rlabel metal1 s 9752 13294 9752 13294 4 _059_
rlabel metal1 s 10718 8262 10718 8262 4 _060_
rlabel metal1 s 11178 8398 11178 8398 4 _061_
rlabel metal1 s 9154 9452 9154 9452 4 _062_
rlabel metal1 s 9384 10574 9384 10574 4 _063_
rlabel metal1 s 7728 9078 7728 9078 4 _064_
rlabel metal1 s 15870 6766 15870 6766 4 _065_
rlabel metal1 s 11132 8330 11132 8330 4 _066_
rlabel metal2 s 10994 8772 10994 8772 4 _067_
rlabel metal1 s 9062 9010 9062 9010 4 _068_
rlabel metal1 s 7774 8806 7774 8806 4 _069_
rlabel metal1 s 9292 8602 9292 8602 4 _070_
rlabel metal1 s 9798 8058 9798 8058 4 _071_
rlabel metal1 s 8786 8432 8786 8432 4 _072_
rlabel metal1 s 3864 7854 3864 7854 4 _073_
rlabel metal1 s 11592 10438 11592 10438 4 _074_
rlabel metal1 s 10212 11322 10212 11322 4 _075_
rlabel metal2 s 9522 10914 9522 10914 4 _076_
rlabel metal1 s 9062 10506 9062 10506 4 _077_
rlabel metal1 s 9798 8296 9798 8296 4 _078_
rlabel metal1 s 7498 7344 7498 7344 4 _079_
rlabel metal1 s 7038 7310 7038 7310 4 _080_
rlabel metal1 s 10350 12614 10350 12614 4 _081_
rlabel metal1 s 15456 8262 15456 8262 4 _082_
rlabel metal2 s 13202 10370 13202 10370 4 _083_
rlabel metal1 s 17204 9010 17204 9010 4 _084_
rlabel metal1 s 15502 10676 15502 10676 4 _085_
rlabel metal1 s 10626 10642 10626 10642 4 _086_
rlabel metal1 s 7866 7276 7866 7276 4 _087_
rlabel metal1 s 6302 7514 6302 7514 4 _088_
rlabel metal2 s 6762 10404 6762 10404 4 _089_
rlabel metal1 s 5336 10438 5336 10438 4 _090_
rlabel metal1 s 7452 6766 7452 6766 4 _091_
rlabel metal1 s 6992 8398 6992 8398 4 _092_
rlabel metal1 s 6954 9078 6954 9078 4 _093_
rlabel metal2 s 7130 9860 7130 9860 4 _094_
rlabel metal1 s 7130 9622 7130 9622 4 _095_
rlabel metal2 s 7222 10132 7222 10132 4 _096_
rlabel metal1 s 14214 10030 14214 10030 4 _097_
rlabel metal1 s 8786 5100 8786 5100 4 _098_
rlabel metal2 s 11178 9894 11178 9894 4 _099_
rlabel metal1 s 11914 10098 11914 10098 4 _100_
rlabel metal1 s 14904 8602 14904 8602 4 _101_
rlabel metal1 s 11914 9010 11914 9010 4 _102_
rlabel metal1 s 13938 11696 13938 11696 4 _103_
rlabel metal1 s 5382 9554 5382 9554 4 _104_
rlabel metal2 s 7498 10404 7498 10404 4 _105_
rlabel metal1 s 6762 10472 6762 10472 4 _106_
rlabel metal1 s 6440 8398 6440 8398 4 _107_
rlabel metal2 s 15225 10098 15225 10098 4 _108_
rlabel metal1 s 5934 6970 5934 6970 4 _109_
rlabel metal1 s 6624 4794 6624 4794 4 _110_
rlabel metal1 s 6808 7718 6808 7718 4 _111_
rlabel metal1 s 8234 4658 8234 4658 4 _112_
rlabel metal2 s 7682 9316 7682 9316 4 _113_
rlabel metal2 s 7682 10438 7682 10438 4 _114_
rlabel metal1 s 6026 8364 6026 8364 4 _115_
rlabel metal1 s 5934 7922 5934 7922 4 _116_
rlabel metal1 s 4784 8330 4784 8330 4 _117_
rlabel metal1 s 5474 8024 5474 8024 4 _118_
rlabel metal1 s 4646 8432 4646 8432 4 _119_
rlabel metal1 s 4094 8058 4094 8058 4 _120_
rlabel metal1 s 4462 8602 4462 8602 4 _121_
rlabel metal1 s 4830 9554 4830 9554 4 _122_
rlabel metal1 s 4738 9486 4738 9486 4 _123_
rlabel metal1 s 4600 9690 4600 9690 4 _124_
rlabel metal1 s 4140 10574 4140 10574 4 _125_
rlabel metal2 s 5842 9044 5842 9044 4 _126_
rlabel metal1 s 6486 9622 6486 9622 4 _127_
rlabel metal1 s 6486 9486 6486 9486 4 _128_
rlabel metal2 s 6394 10098 6394 10098 4 _129_
rlabel metal1 s 4094 7310 4094 7310 4 _130_
rlabel metal1 s 4876 7990 4876 7990 4 _131_
rlabel metal1 s 4922 7888 4922 7888 4 _132_
rlabel metal1 s 4140 7514 4140 7514 4 _133_
rlabel metal2 s 5106 6426 5106 6426 4 _134_
rlabel metal1 s 5014 6086 5014 6086 4 _135_
rlabel metal1 s 3818 6426 3818 6426 4 _136_
rlabel metal1 s 3818 7310 3818 7310 4 _137_
rlabel metal1 s 6440 5270 6440 5270 4 _138_
rlabel metal2 s 5658 5984 5658 5984 4 _139_
rlabel metal1 s 5198 5780 5198 5780 4 _140_
rlabel metal2 s 5842 5270 5842 5270 4 _141_
rlabel metal1 s 6440 5202 6440 5202 4 _142_
rlabel metal1 s 7452 6222 7452 6222 4 _143_
rlabel metal1 s 6854 5814 6854 5814 4 _144_
rlabel metal1 s 7314 4726 7314 4726 4 _145_
rlabel metal1 s 6348 5338 6348 5338 4 _146_
rlabel metal1 s 7406 5134 7406 5134 4 _147_
rlabel metal2 s 7958 4828 7958 4828 4 _148_
rlabel metal2 s 7866 4607 7866 4607 4 _149_
rlabel metal1 s 7912 4522 7912 4522 4 _150_
rlabel metal2 s 8694 4352 8694 4352 4 _151_
rlabel metal1 s 9844 3570 9844 3570 4 _152_
rlabel metal2 s 13110 13838 13110 13838 4 _153_
rlabel metal1 s 6624 13430 6624 13430 4 _154_
rlabel metal1 s 2714 13226 2714 13226 4 _155_
rlabel metal2 s 8142 17510 8142 17510 4 _156_
rlabel metal1 s 7682 16048 7682 16048 4 _157_
rlabel metal1 s 6348 17578 6348 17578 4 _158_
rlabel metal1 s 6486 17510 6486 17510 4 _159_
rlabel metal1 s 6440 17850 6440 17850 4 _160_
rlabel metal2 s 5566 16286 5566 16286 4 _161_
rlabel metal2 s 4738 17816 4738 17816 4 _162_
rlabel metal1 s 4508 17714 4508 17714 4 _163_
rlabel metal1 s 5152 16150 5152 16150 4 _164_
rlabel metal1 s 5060 16218 5060 16218 4 _165_
rlabel metal1 s 4646 16014 4646 16014 4 _166_
rlabel metal2 s 6394 15164 6394 15164 4 _167_
rlabel metal2 s 6026 14790 6026 14790 4 _168_
rlabel metal1 s 5290 14586 5290 14586 4 _169_
rlabel metal2 s 6210 13600 6210 13600 4 _170_
rlabel metal2 s 6578 13430 6578 13430 4 _171_
rlabel metal1 s 6946 13226 6946 13226 4 _172_
rlabel metal2 s 5842 12517 5842 12517 4 _173_
rlabel metal1 s 4646 13362 4646 13362 4 _174_
rlabel metal1 s 4784 13498 4784 13498 4 _175_
rlabel metal1 s 4646 12274 4646 12274 4 _176_
rlabel metal2 s 3266 14144 3266 14144 4 _177_
rlabel metal1 s 2438 13396 2438 13396 4 _178_
rlabel metal1 s 4002 14280 4002 14280 4 _179_
rlabel metal1 s 4132 14586 4132 14586 4 _180_
rlabel metal1 s 2530 13872 2530 13872 4 _181_
rlabel metal2 s 3450 15164 3450 15164 4 _182_
rlabel metal1 s 3174 14926 3174 14926 4 _183_
rlabel metal1 s 11546 14858 11546 14858 4 _184_
rlabel metal2 s 13754 13583 13754 13583 4 _185_
rlabel metal2 s 13662 13532 13662 13532 4 _186_
rlabel metal1 s 12880 13702 12880 13702 4 _187_
rlabel metal2 s 13110 4862 13110 4862 4 _188_
rlabel metal1 s 13202 7311 13202 7311 4 _189_
rlabel metal2 s 13570 5372 13570 5372 4 _190_
rlabel metal1 s 13110 8976 13110 8976 4 _191_
rlabel metal2 s 13478 6188 13478 6188 4 _192_
rlabel metal2 s 12834 7140 12834 7140 4 _193_
rlabel metal2 s 12742 7412 12742 7412 4 _194_
rlabel metal1 s 12696 7990 12696 7990 4 _195_
rlabel metal1 s 12834 9554 12834 9554 4 _196_
rlabel metal1 s 12144 9690 12144 9690 4 _197_
rlabel metal2 s 16790 8602 16790 8602 4 _198_
rlabel metal2 s 16146 5440 16146 5440 4 _199_
rlabel metal1 s 15962 9418 15962 9418 4 _200_
rlabel metal1 s 14996 9690 14996 9690 4 _201_
rlabel metal1 s 15042 10064 15042 10064 4 _202_
rlabel metal1 s 12466 10030 12466 10030 4 _203_
rlabel metal1 s 12052 10234 12052 10234 4 _204_
rlabel metal2 s 11914 11764 11914 11764 4 _205_
rlabel metal1 s 11316 12274 11316 12274 4 _206_
rlabel metal1 s 13432 12682 13432 12682 4 _207_
rlabel metal1 s 15847 9486 15847 9486 4 _208_
rlabel metal1 s 16008 10574 16008 10574 4 _209_
rlabel metal1 s 15502 9520 15502 9520 4 _210_
rlabel metal2 s 15870 10438 15870 10438 4 _211_
rlabel metal2 s 13754 9010 13754 9010 4 _212_
rlabel metal2 s 14043 9486 14043 9486 4 _213_
rlabel metal1 s 13984 9146 13984 9146 4 _214_
rlabel metal1 s 13432 9690 13432 9690 4 _215_
rlabel metal1 s 13478 9350 13478 9350 4 _216_
rlabel metal1 s 13570 10234 13570 10234 4 _217_
rlabel metal2 s 14030 11730 14030 11730 4 _218_
rlabel metal1 s 13616 12750 13616 12750 4 _219_
rlabel metal2 s 12374 12818 12374 12818 4 _220_
rlabel metal1 s 16697 7922 16697 7922 4 _221_
rlabel metal1 s 16606 7344 16606 7344 4 _222_
rlabel metal2 s 15410 7344 15410 7344 4 _223_
rlabel metal2 s 15502 5508 15502 5508 4 _224_
rlabel metal2 s 15962 6562 15962 6562 4 _225_
rlabel metal1 s 16468 6834 16468 6834 4 _226_
rlabel metal1 s 16514 6188 16514 6188 4 _227_
rlabel metal1 s 17204 6086 17204 6086 4 _228_
rlabel metal2 s 16330 7174 16330 7174 4 _229_
rlabel metal1 s 16422 7514 16422 7514 4 _230_
rlabel metal1 s 15502 7888 15502 7888 4 _231_
rlabel metal1 s 14490 8058 14490 8058 4 _232_
rlabel metal1 s 14858 8432 14858 8432 4 _233_
rlabel metal1 s 13846 8432 13846 8432 4 _234_
rlabel metal1 s 13754 8466 13754 8466 4 _235_
rlabel metal2 s 13570 10404 13570 10404 4 _236_
rlabel metal1 s 12742 12410 12742 12410 4 _237_
rlabel metal3 s 10327 18020 10327 18020 4 _238_
rlabel metal1 s 14582 5236 14582 5236 4 _239_
rlabel metal2 s 14674 5270 14674 5270 4 _240_
rlabel metal2 s 14214 5610 14214 5610 4 _241_
rlabel metal2 s 14122 4828 14122 4828 4 _242_
rlabel metal2 s 14950 5372 14950 5372 4 _243_
rlabel metal1 s 13754 5338 13754 5338 4 _244_
rlabel metal2 s 15686 6630 15686 6630 4 _245_
rlabel metal2 s 14674 6494 14674 6494 4 _246_
rlabel metal2 s 15042 6018 15042 6018 4 _247_
rlabel metal1 s 13386 5780 13386 5780 4 _248_
rlabel metal1 s 12696 5882 12696 5882 4 _249_
rlabel metal1 s 11132 11866 11132 11866 4 _250_
rlabel metal1 s 10580 12614 10580 12614 4 _251_
rlabel metal1 s 15410 4726 15410 4726 4 _252_
rlabel metal1 s 14858 4046 14858 4046 4 _253_
rlabel metal2 s 14582 4454 14582 4454 4 _254_
rlabel metal1 s 14674 4794 14674 4794 4 _255_
rlabel metal2 s 12742 4964 12742 4964 4 _256_
rlabel metal2 s 12466 4964 12466 4964 4 _257_
rlabel metal3 s 12926 5355 12926 5355 4 _258_
rlabel metal1 s 11868 12410 11868 12410 4 _259_
rlabel metal2 s 11546 14008 11546 14008 4 _260_
rlabel metal1 s 14260 4250 14260 4250 4 _261_
rlabel metal1 s 12558 4012 12558 4012 4 _262_
rlabel metal1 s 11868 13974 11868 13974 4 _263_
rlabel metal1 s 11684 13838 11684 13838 4 _264_
rlabel metal1 s 11868 12614 11868 12614 4 _265_
rlabel metal1 s 12604 7310 12604 7310 4 _266_
rlabel metal1 s 12144 6970 12144 6970 4 _267_
rlabel metal1 s 13018 13906 13018 13906 4 _268_
rlabel metal2 s 12558 13260 12558 13260 4 _269_
rlabel metal1 s 13248 11866 13248 11866 4 _270_
rlabel metal1 s 13662 13906 13662 13906 4 _271_
rlabel metal2 s 14398 11356 14398 11356 4 _272_
rlabel metal1 s 13708 14042 13708 14042 4 _273_
rlabel metal1 s 13202 17680 13202 17680 4 _274_
rlabel metal2 s 15594 10387 15594 10387 4 _275_
rlabel metal1 s 8694 16558 8694 16558 4 _276_
rlabel metal1 s 9155 15504 9155 15504 4 _277_
rlabel metal1 s 8924 16014 8924 16014 4 _278_
rlabel metal1 s 10028 8466 10028 8466 4 _279_
rlabel metal1 s 7774 14416 7774 14416 4 _280_
rlabel metal2 s 7958 14246 7958 14246 4 _281_
rlabel metal1 s 7958 14518 7958 14518 4 _282_
rlabel metal2 s 19090 14613 19090 14613 4 clk
rlabel metal1 s 10028 13430 10028 13430 4 clknet_0_clk
rlabel metal1 s 4922 4046 4922 4046 4 clknet_2_0__leaf_clk
rlabel metal1 s 13294 1360 13294 1360 4 clknet_2_1__leaf_clk
rlabel metal1 s 6026 18190 6026 18190 4 clknet_2_2__leaf_clk
rlabel metal1 s 12466 16592 12466 16592 4 clknet_2_3__leaf_clk
rlabel metal1 s 16054 18802 16054 18802 4 data[0]
rlabel metal1 s 14260 18802 14260 18802 4 data[1]
rlabel metal1 s 12512 18802 12512 18802 4 data[2]
rlabel metal1 s 10994 18802 10994 18802 4 data[3]
rlabel metal1 s 9200 18802 9200 18802 4 data[4]
rlabel metal1 s 7544 18802 7544 18802 4 data[5]
rlabel metal1 s 5888 18802 5888 18802 4 data[6]
rlabel metal1 s 4232 18802 4232 18802 4 data[7]
rlabel metal1 s 2576 18802 2576 18802 4 ext_data
rlabel metal1 s 920 18802 920 18802 4 load_divider
rlabel metal1 s 17572 18802 17572 18802 4 n_rst
rlabel metal2 s 16146 17408 16146 17408 4 net1
rlabel metal1 s 7682 15640 7682 15640 4 net10
rlabel metal2 s 16698 18394 16698 18394 4 net11
rlabel metal2 s 15134 17408 15134 17408 4 net12
rlabel metal1 s 8556 14518 8556 14518 4 net13
rlabel metal1 s 10718 17782 10718 17782 4 net14
rlabel metal1 s 7912 15606 7912 15606 4 net15
rlabel metal1 s 10304 16694 10304 16694 4 net16
rlabel metal1 s 10304 15606 10304 15606 4 net17
rlabel metal1 s 12788 17782 12788 17782 4 net18
rlabel metal1 s 11914 17000 11914 17000 4 net19
rlabel metal2 s 13570 17306 13570 17306 4 net2
rlabel metal2 s 11546 15810 11546 15810 4 net20
rlabel metal1 s 3220 13294 3220 13294 4 net21
rlabel metal2 s 7866 16320 7866 16320 4 net22
rlabel metal1 s 6670 16218 6670 16218 4 net23
rlabel metal1 s 13938 13872 13938 13872 4 net24
rlabel metal1 s 6164 12614 6164 12614 4 net25
rlabel metal1 s 12788 18598 12788 18598 4 net3
rlabel metal2 s 10350 18394 10350 18394 4 net4
rlabel metal2 s 10350 16847 10350 16847 4 net5
rlabel metal1 s 7590 15504 7590 15504 4 net6
rlabel metal1 s 10442 15538 10442 15538 4 net7
rlabel metal2 s 13938 13804 13938 13804 4 net8
rlabel metal2 s 12558 16830 12558 16830 4 net9
rlabel metal2 s 1242 942 1242 942 4 r2r_out[0]
rlabel metal2 s 12834 2720 12834 2720 4 r2r_out[1]
rlabel metal1 s 9016 2822 9016 2822 4 r2r_out[2]
rlabel metal2 s 8694 1486 8694 1486 4 r2r_out[3]
rlabel metal2 s 11178 1044 11178 1044 4 r2r_out[4]
rlabel metal2 s 13662 942 13662 942 4 r2r_out[5]
rlabel metal2 s 16146 500 16146 500 4 r2r_out[6]
rlabel metal2 s 18630 942 18630 942 4 r2r_out[7]
rlabel metal1 s 9614 16728 9614 16728 4 sine_lookup.count\[0\]
rlabel metal1 s 3542 14552 3542 14552 4 sine_lookup.count\[10\]
rlabel metal1 s 4278 15538 4278 15538 4 sine_lookup.count\[11\]
rlabel metal1 s 7406 17544 7406 17544 4 sine_lookup.count\[1\]
rlabel metal1 s 7222 18292 7222 18292 4 sine_lookup.count\[2\]
rlabel metal1 s 6256 17646 6256 17646 4 sine_lookup.count\[3\]
rlabel metal1 s 6118 15946 6118 15946 4 sine_lookup.count\[4\]
rlabel metal2 s 6026 15912 6026 15912 4 sine_lookup.count\[5\]
rlabel metal1 s 8372 13838 8372 13838 4 sine_lookup.count\[6\]
rlabel metal1 s 7590 13804 7590 13804 4 sine_lookup.count\[7\]
rlabel metal1 s 5198 14008 5198 14008 4 sine_lookup.count\[8\]
rlabel metal1 s 4232 13838 4232 13838 4 sine_lookup.count\[9\]
rlabel metal2 s 13110 15708 13110 15708 4 sine_lookup.divider\[0\]
rlabel metal2 s 13018 16932 13018 16932 4 sine_lookup.divider\[1\]
rlabel metal1 s 9890 18394 9890 18394 4 sine_lookup.divider\[2\]
rlabel metal1 s 10074 18326 10074 18326 4 sine_lookup.divider\[3\]
rlabel metal2 s 10994 16286 10994 16286 4 sine_lookup.divider\[4\]
rlabel metal1 s 7774 14790 7774 14790 4 sine_lookup.divider\[5\]
rlabel metal2 s 10994 15844 10994 15844 4 sine_lookup.divider\[6\]
rlabel metal2 s 9430 14212 9430 14212 4 sine_lookup.divider\[7\]
rlabel metal1 s 9591 8466 9591 8466 4 sine_lookup.rst
rlabel metal1 s 11178 10506 11178 10506 4 sine_lookup.sine_input\[0\]
rlabel metal1 s 15042 8364 15042 8364 4 sine_lookup.sine_input\[1\]
rlabel metal1 s 10212 6698 10212 6698 4 sine_lookup.sine_input\[2\]
rlabel metal2 s 10534 6783 10534 6783 4 sine_lookup.sine_input\[3\]
rlabel metal2 s 12650 7310 12650 7310 4 sine_lookup.sine_input\[4\]
rlabel metal1 s 13478 10132 13478 10132 4 sine_lookup.sine_input\[5\]
rlabel metal1 s 13432 5134 13432 5134 4 sine_lookup.sine_input\[6\]
rlabel metal1 s 15042 14348 15042 14348 4 sine_lookup.sine_input\[7\]
flabel metal4 s 19251 496 19571 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14536 496 14856 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9821 496 10141 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5106 496 5426 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16894 496 17214 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12179 496 12499 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7464 496 7784 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2749 496 3069 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 19062 19600 19118 20000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 15750 19600 15806 20000 0 FreeSans 280 90 0 0 data[0]
port 4 nsew
flabel metal2 s 14094 19600 14150 20000 0 FreeSans 280 90 0 0 data[1]
port 5 nsew
flabel metal2 s 12438 19600 12494 20000 0 FreeSans 280 90 0 0 data[2]
port 6 nsew
flabel metal2 s 10782 19600 10838 20000 0 FreeSans 280 90 0 0 data[3]
port 7 nsew
flabel metal2 s 9126 19600 9182 20000 0 FreeSans 280 90 0 0 data[4]
port 8 nsew
flabel metal2 s 7470 19600 7526 20000 0 FreeSans 280 90 0 0 data[5]
port 9 nsew
flabel metal2 s 5814 19600 5870 20000 0 FreeSans 280 90 0 0 data[6]
port 10 nsew
flabel metal2 s 4158 19600 4214 20000 0 FreeSans 280 90 0 0 data[7]
port 11 nsew
flabel metal2 s 2502 19600 2558 20000 0 FreeSans 280 90 0 0 ext_data
port 12 nsew
flabel metal2 s 846 19600 902 20000 0 FreeSans 280 90 0 0 load_divider
port 13 nsew
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 280 90 0 0 n_rst
port 14 nsew
flabel metal2 s 1214 0 1270 400 0 FreeSans 280 90 0 0 r2r_out[0]
port 15 nsew
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 r2r_out[1]
port 16 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 r2r_out[2]
port 17 nsew
flabel metal2 s 8666 0 8722 400 0 FreeSans 280 90 0 0 r2r_out[3]
port 18 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 r2r_out[4]
port 19 nsew
flabel metal2 s 13634 0 13690 400 0 FreeSans 280 90 0 0 r2r_out[5]
port 20 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 r2r_out[6]
port 21 nsew
flabel metal2 s 18602 0 18658 400 0 FreeSans 280 90 0 0 r2r_out[7]
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string GDS_END 1359276
string GDS_FILE ../gds/r2r_dac_control.gds
string GDS_START 395382
<< end >>
