magic
tech sky130A
magscale 1 2
timestamp 1720092317
<< nwell >>
rect -308 -346 308 346
<< mvpmos >>
rect -50 -120 50 48
<< mvpdiff >>
rect -108 36 -50 48
rect -108 -108 -96 36
rect -62 -108 -50 36
rect -108 -120 -50 -108
rect 50 36 108 48
rect 50 -108 62 36
rect 96 -108 108 36
rect 50 -120 108 -108
<< mvpdiffc >>
rect -96 -108 -62 36
rect 62 -108 96 36
<< mvnsubdiff >>
rect -242 268 242 280
rect -242 234 -134 268
rect 134 234 242 268
rect -242 222 242 234
rect -242 172 -184 222
rect -242 -172 -230 172
rect -196 -172 -184 172
rect 184 172 242 222
rect -242 -222 -184 -172
rect 184 -172 196 172
rect 230 -172 242 172
rect 184 -222 242 -172
rect -242 -234 242 -222
rect -242 -268 -134 -234
rect 134 -268 242 -234
rect -242 -280 242 -268
<< mvnsubdiffcont >>
rect -134 234 134 268
rect -230 -172 -196 172
rect 196 -172 230 172
rect -134 -268 134 -234
<< poly >>
rect -50 129 50 145
rect -50 95 -34 129
rect 34 95 50 129
rect -50 48 50 95
rect -50 -146 50 -120
<< polycont >>
rect -34 95 34 129
<< locali >>
rect -230 234 -134 268
rect 134 234 230 268
rect -230 172 -196 234
rect 196 172 230 234
rect -50 95 -34 129
rect 34 95 50 129
rect -96 36 -62 52
rect -96 -124 -62 -108
rect 62 36 96 52
rect 62 -124 96 -108
rect -230 -234 -196 -172
rect 196 -234 230 -172
rect -230 -268 -134 -234
rect 134 -268 230 -234
<< viali >>
rect -34 95 34 129
rect -96 -108 -62 36
rect 62 -108 96 36
<< metal1 >>
rect -46 129 46 135
rect -46 95 -34 129
rect 34 95 46 129
rect -46 89 46 95
rect -102 36 -56 48
rect -102 -108 -96 36
rect -62 -108 -56 36
rect -102 -120 -56 -108
rect 56 36 102 48
rect 56 -108 62 36
rect 96 -108 102 36
rect 56 -120 102 -108
<< properties >>
string FIXED_BBOX -213 -251 213 251
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.84 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
