magic
tech sky130A
magscale 1 2
timestamp 1720104585
<< viali >>
rect 949 18785 983 18819
rect 2605 18785 2639 18819
rect 4261 18785 4295 18819
rect 5917 18785 5951 18819
rect 7573 18785 7607 18819
rect 8953 18785 8987 18819
rect 9597 18785 9631 18819
rect 10977 18785 11011 18819
rect 12725 18785 12759 18819
rect 14381 18785 14415 18819
rect 16313 18785 16347 18819
rect 17693 18785 17727 18819
rect 1225 18717 1259 18751
rect 8861 18717 8895 18751
rect 9321 18717 9355 18751
rect 2789 18649 2823 18683
rect 16129 18649 16163 18683
rect 4445 18581 4479 18615
rect 6101 18581 6135 18615
rect 7757 18581 7791 18615
rect 8677 18581 8711 18615
rect 9413 18581 9447 18615
rect 11161 18581 11195 18615
rect 12541 18581 12575 18615
rect 14197 18581 14231 18615
rect 17509 18581 17543 18615
rect 7113 18377 7147 18411
rect 6837 18309 6871 18343
rect 9781 18309 9815 18343
rect 5457 18173 5491 18207
rect 6929 18173 6963 18207
rect 7297 18173 7331 18207
rect 8401 18173 8435 18207
rect 8668 18173 8702 18207
rect 9873 18173 9907 18207
rect 11069 18173 11103 18207
rect 13093 18173 13127 18207
rect 13185 18173 13219 18207
rect 14933 18173 14967 18207
rect 15117 18173 15151 18207
rect 17141 18173 17175 18207
rect 5724 18105 5758 18139
rect 11336 18105 11370 18139
rect 13369 18105 13403 18139
rect 14666 18105 14700 18139
rect 15393 18105 15427 18139
rect 17049 18105 17083 18139
rect 7389 18037 7423 18071
rect 9965 18037 9999 18071
rect 12449 18037 12483 18071
rect 12725 18037 12759 18071
rect 13553 18037 13587 18071
rect 16865 18037 16899 18071
rect 6009 17833 6043 17867
rect 6653 17833 6687 17867
rect 6745 17833 6779 17867
rect 8861 17833 8895 17867
rect 12357 17833 12391 17867
rect 13001 17833 13035 17867
rect 15485 17833 15519 17867
rect 6285 17697 6319 17731
rect 6929 17697 6963 17731
rect 7113 17697 7147 17731
rect 7656 17697 7690 17731
rect 9229 17697 9263 17731
rect 9413 17697 9447 17731
rect 9680 17697 9714 17731
rect 10977 17697 11011 17731
rect 11253 17697 11287 17731
rect 12081 17697 12115 17731
rect 12449 17697 12483 17731
rect 13277 17697 13311 17731
rect 13369 17697 13403 17731
rect 13645 17697 13679 17731
rect 13737 17697 13771 17731
rect 6193 17629 6227 17663
rect 7389 17629 7423 17663
rect 9137 17629 9171 17663
rect 11161 17629 11195 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 12173 17629 12207 17663
rect 7113 17493 7147 17527
rect 8769 17493 8803 17527
rect 9229 17493 9263 17527
rect 10793 17493 10827 17527
rect 12541 17493 12575 17527
rect 13369 17493 13403 17527
rect 13553 17493 13587 17527
rect 13829 17493 13863 17527
rect 7205 17289 7239 17323
rect 8033 17289 8067 17323
rect 9045 17289 9079 17323
rect 10333 17289 10367 17323
rect 10517 17289 10551 17323
rect 10977 17289 11011 17323
rect 11253 17289 11287 17323
rect 6469 17153 6503 17187
rect 7941 17153 7975 17187
rect 8861 17153 8895 17187
rect 10241 17153 10275 17187
rect 10977 17153 11011 17187
rect 13553 17153 13587 17187
rect 4813 17085 4847 17119
rect 6561 17085 6595 17119
rect 7205 17085 7239 17119
rect 7389 17085 7423 17119
rect 7849 17085 7883 17119
rect 8769 17085 8803 17119
rect 9137 17085 9171 17119
rect 10149 17085 10183 17119
rect 10885 17085 10919 17119
rect 11529 17085 11563 17119
rect 11621 17085 11655 17119
rect 12173 17085 12207 17119
rect 13093 17085 13127 17119
rect 13185 17085 13219 17119
rect 5080 17017 5114 17051
rect 6285 17017 6319 17051
rect 11713 17017 11747 17051
rect 13369 17017 13403 17051
rect 13798 17017 13832 17051
rect 6193 16949 6227 16983
rect 6929 16949 6963 16983
rect 7021 16949 7055 16983
rect 8217 16949 8251 16983
rect 8401 16949 8435 16983
rect 9229 16949 9263 16983
rect 11437 16949 11471 16983
rect 12357 16949 12391 16983
rect 12725 16949 12759 16983
rect 14933 16949 14967 16983
rect 9321 16745 9355 16779
rect 12909 16745 12943 16779
rect 6469 16677 6503 16711
rect 6377 16609 6411 16643
rect 6653 16609 6687 16643
rect 6929 16609 6963 16643
rect 7021 16609 7055 16643
rect 8677 16609 8711 16643
rect 9229 16609 9263 16643
rect 13277 16609 13311 16643
rect 13921 16609 13955 16643
rect 6745 16541 6779 16575
rect 13185 16541 13219 16575
rect 7205 16405 7239 16439
rect 8861 16405 8895 16439
rect 9137 16405 9171 16439
rect 13277 16405 13311 16439
rect 13829 16405 13863 16439
rect 6469 16133 6503 16167
rect 7297 16133 7331 16167
rect 9413 16133 9447 16167
rect 12817 16065 12851 16099
rect 12909 16065 12943 16099
rect 6193 15997 6227 16031
rect 6285 15997 6319 16031
rect 6653 15997 6687 16031
rect 6801 15997 6835 16031
rect 7021 15997 7055 16031
rect 7159 15997 7193 16031
rect 7573 15997 7607 16031
rect 7757 15997 7791 16031
rect 7941 15997 7975 16031
rect 8769 15997 8803 16031
rect 8861 15997 8895 16031
rect 9229 15997 9263 16031
rect 9505 15997 9539 16031
rect 9689 15997 9723 16031
rect 9781 15997 9815 16031
rect 9873 15997 9907 16031
rect 10057 15997 10091 16031
rect 10977 15997 11011 16031
rect 11069 15997 11103 16031
rect 11161 15997 11195 16031
rect 11345 15997 11379 16031
rect 12633 15997 12667 16031
rect 13001 15997 13035 16031
rect 13185 15997 13219 16031
rect 13553 15997 13587 16031
rect 13737 15997 13771 16031
rect 13829 15997 13863 16031
rect 14013 15997 14047 16031
rect 14105 15997 14139 16031
rect 6929 15929 6963 15963
rect 7665 15929 7699 15963
rect 9045 15929 9079 15963
rect 9137 15929 9171 15963
rect 6101 15861 6135 15895
rect 7389 15861 7423 15895
rect 10241 15861 10275 15895
rect 10793 15861 10827 15895
rect 12449 15861 12483 15895
rect 6469 15657 6503 15691
rect 7849 15657 7883 15691
rect 9137 15657 9171 15691
rect 14197 15657 14231 15691
rect 7389 15589 7423 15623
rect 8861 15589 8895 15623
rect 9597 15589 9631 15623
rect 4528 15521 4562 15555
rect 6653 15521 6687 15555
rect 6929 15521 6963 15555
rect 7113 15521 7147 15555
rect 8585 15521 8619 15555
rect 8769 15521 8803 15555
rect 8953 15521 8987 15555
rect 10149 15521 10183 15555
rect 10333 15521 10367 15555
rect 10425 15521 10459 15555
rect 10517 15521 10551 15555
rect 11233 15521 11267 15555
rect 12909 15521 12943 15555
rect 4261 15453 4295 15487
rect 10057 15453 10091 15487
rect 10977 15453 11011 15487
rect 7665 15385 7699 15419
rect 9965 15385 9999 15419
rect 5641 15317 5675 15351
rect 10793 15317 10827 15351
rect 12357 15317 12391 15351
rect 5089 15113 5123 15147
rect 10701 15113 10735 15147
rect 12357 15113 12391 15147
rect 13553 15113 13587 15147
rect 6745 15045 6779 15079
rect 7665 14977 7699 15011
rect 14933 14977 14967 15011
rect 5273 14909 5307 14943
rect 6285 14909 6319 14943
rect 6469 14909 6503 14943
rect 6561 14909 6595 14943
rect 7389 14909 7423 14943
rect 7481 14909 7515 14943
rect 10517 14909 10551 14943
rect 12817 14909 12851 14943
rect 6929 14841 6963 14875
rect 12173 14841 12207 14875
rect 14666 14841 14700 14875
rect 6101 14773 6135 14807
rect 7021 14773 7055 14807
rect 7113 14773 7147 14807
rect 7297 14773 7331 14807
rect 7665 14773 7699 14807
rect 12373 14773 12407 14807
rect 12541 14773 12575 14807
rect 13001 14773 13035 14807
rect 10333 14569 10367 14603
rect 10425 14569 10459 14603
rect 11345 14569 11379 14603
rect 12265 14569 12299 14603
rect 5441 14501 5475 14535
rect 5641 14501 5675 14535
rect 6561 14501 6595 14535
rect 9029 14501 9063 14535
rect 9229 14501 9263 14535
rect 9781 14501 9815 14535
rect 10577 14501 10611 14535
rect 10793 14501 10827 14535
rect 11713 14501 11747 14535
rect 11805 14501 11839 14535
rect 12633 14501 12667 14535
rect 12985 14501 13019 14535
rect 13185 14501 13219 14535
rect 6193 14433 6227 14467
rect 6285 14433 6319 14467
rect 8769 14433 8803 14467
rect 10057 14433 10091 14467
rect 11161 14433 11195 14467
rect 11437 14433 11471 14467
rect 11897 14433 11931 14467
rect 12449 14433 12483 14467
rect 12725 14433 12759 14467
rect 6653 14365 6687 14399
rect 7021 14365 7055 14399
rect 9689 14365 9723 14399
rect 10149 14365 10183 14399
rect 5273 14297 5307 14331
rect 6009 14297 6043 14331
rect 8861 14297 8895 14331
rect 12081 14297 12115 14331
rect 12817 14297 12851 14331
rect 5457 14229 5491 14263
rect 9045 14229 9079 14263
rect 10609 14229 10643 14263
rect 10977 14229 11011 14263
rect 11529 14229 11563 14263
rect 13001 14229 13035 14263
rect 6837 14025 6871 14059
rect 8401 14025 8435 14059
rect 12357 14025 12391 14059
rect 5733 13957 5767 13991
rect 13553 13957 13587 13991
rect 6377 13889 6411 13923
rect 6469 13889 6503 13923
rect 8217 13889 8251 13923
rect 9597 13889 9631 13923
rect 11805 13889 11839 13923
rect 12817 13889 12851 13923
rect 14933 13889 14967 13923
rect 4353 13821 4387 13855
rect 4620 13821 4654 13855
rect 6009 13821 6043 13855
rect 6193 13821 6227 13855
rect 6561 13821 6595 13855
rect 6745 13821 6779 13855
rect 8401 13821 8435 13855
rect 8585 13821 8619 13855
rect 8953 13821 8987 13855
rect 9137 13821 9171 13855
rect 9229 13821 9263 13855
rect 9321 13821 9355 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 12081 13821 12115 13855
rect 12173 13821 12207 13855
rect 12449 13821 12483 13855
rect 12633 13821 12667 13855
rect 12725 13821 12759 13855
rect 13001 13821 13035 13855
rect 13185 13821 13219 13855
rect 14666 13821 14700 13855
rect 7950 13753 7984 13787
rect 9689 13753 9723 13787
rect 11713 13753 11747 13787
rect 6009 13481 6043 13515
rect 7665 13481 7699 13515
rect 7849 13481 7883 13515
rect 8795 13481 8829 13515
rect 12725 13481 12759 13515
rect 13001 13481 13035 13515
rect 8585 13413 8619 13447
rect 10158 13413 10192 13447
rect 6193 13345 6227 13379
rect 6929 13345 6963 13379
rect 7113 13345 7147 13379
rect 7205 13345 7239 13379
rect 7481 13345 7515 13379
rect 7757 13345 7791 13379
rect 7941 13345 7975 13379
rect 10425 13345 10459 13379
rect 12541 13345 12575 13379
rect 12817 13345 12851 13379
rect 13093 13345 13127 13379
rect 6377 13277 6411 13311
rect 7297 13277 7331 13311
rect 12357 13277 12391 13311
rect 9045 13209 9079 13243
rect 12817 13209 12851 13243
rect 8769 13141 8803 13175
rect 8953 13141 8987 13175
rect 6653 12937 6687 12971
rect 9137 12937 9171 12971
rect 11529 12937 11563 12971
rect 14933 12937 14967 12971
rect 10057 12869 10091 12903
rect 5733 12801 5767 12835
rect 9689 12801 9723 12835
rect 11805 12801 11839 12835
rect 12173 12801 12207 12835
rect 12633 12801 12667 12835
rect 5273 12733 5307 12767
rect 5365 12733 5399 12767
rect 5457 12733 5491 12767
rect 5641 12733 5675 12767
rect 6377 12733 6411 12767
rect 9321 12733 9355 12767
rect 9413 12733 9447 12767
rect 9873 12733 9907 12767
rect 11345 12733 11379 12767
rect 11989 12733 12023 12767
rect 12265 12733 12299 12767
rect 12449 12733 12483 12767
rect 12541 12733 12575 12767
rect 12817 12733 12851 12767
rect 13553 12733 13587 12767
rect 6469 12665 6503 12699
rect 9781 12665 9815 12699
rect 13001 12665 13035 12699
rect 13798 12665 13832 12699
rect 4997 12597 5031 12631
rect 6669 12597 6703 12631
rect 6837 12597 6871 12631
rect 5917 12393 5951 12427
rect 7205 12393 7239 12427
rect 10149 12393 10183 12427
rect 13001 12393 13035 12427
rect 4436 12325 4470 12359
rect 6929 12325 6963 12359
rect 7021 12325 7055 12359
rect 12725 12325 12759 12359
rect 4169 12257 4203 12291
rect 6193 12257 6227 12291
rect 6837 12257 6871 12291
rect 7573 12257 7607 12291
rect 7757 12257 7791 12291
rect 7849 12257 7883 12291
rect 10333 12257 10367 12291
rect 11069 12257 11103 12291
rect 12817 12257 12851 12291
rect 13093 12257 13127 12291
rect 6101 12189 6135 12223
rect 6469 12189 6503 12223
rect 6561 12189 6595 12223
rect 9689 12189 9723 12223
rect 9781 12189 9815 12223
rect 5549 12121 5583 12155
rect 6653 12121 6687 12155
rect 10517 12121 10551 12155
rect 12817 12121 12851 12155
rect 7573 12053 7607 12087
rect 9505 12053 9539 12087
rect 8033 11849 8067 11883
rect 8125 11849 8159 11883
rect 8401 11849 8435 11883
rect 5457 11781 5491 11815
rect 6377 11713 6411 11747
rect 7297 11713 7331 11747
rect 7665 11713 7699 11747
rect 7941 11713 7975 11747
rect 8861 11713 8895 11747
rect 8953 11713 8987 11747
rect 9873 11713 9907 11747
rect 11529 11713 11563 11747
rect 11713 11713 11747 11747
rect 12265 11713 12299 11747
rect 4077 11645 4111 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 7481 11645 7515 11679
rect 8217 11645 8251 11679
rect 9413 11645 9447 11679
rect 9597 11645 9631 11679
rect 11437 11645 11471 11679
rect 11897 11645 11931 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 12449 11645 12483 11679
rect 13737 11645 13771 11679
rect 4344 11577 4378 11611
rect 7113 11577 7147 11611
rect 7205 11577 7239 11611
rect 9965 11577 9999 11611
rect 12633 11577 12667 11611
rect 5825 11509 5859 11543
rect 6561 11509 6595 11543
rect 8769 11509 8803 11543
rect 9597 11509 9631 11543
rect 10057 11509 10091 11543
rect 10425 11509 10459 11543
rect 11069 11509 11103 11543
rect 13921 11509 13955 11543
rect 5825 11305 5859 11339
rect 10793 11305 10827 11339
rect 12081 11305 12115 11339
rect 13001 11305 13035 11339
rect 10241 11237 10275 11271
rect 13277 11237 13311 11271
rect 6101 11169 6135 11203
rect 6193 11169 6227 11203
rect 6285 11169 6319 11203
rect 6469 11169 6503 11203
rect 7665 11169 7699 11203
rect 10517 11169 10551 11203
rect 11529 11169 11563 11203
rect 11989 11169 12023 11203
rect 12173 11169 12207 11203
rect 12817 11169 12851 11203
rect 7389 11101 7423 11135
rect 8769 11101 8803 11135
rect 10149 11101 10183 11135
rect 10609 11101 10643 11135
rect 11437 11101 11471 11135
rect 12633 11101 12667 11135
rect 11897 11033 11931 11067
rect 14565 10965 14599 10999
rect 10885 10761 10919 10795
rect 11069 10761 11103 10795
rect 7297 10693 7331 10727
rect 10517 10625 10551 10659
rect 10977 10625 11011 10659
rect 13829 10625 13863 10659
rect 7021 10557 7055 10591
rect 7297 10557 7331 10591
rect 7941 10557 7975 10591
rect 10701 10557 10735 10591
rect 11161 10557 11195 10591
rect 11253 10557 11287 10591
rect 11529 10557 11563 10591
rect 13553 10557 13587 10591
rect 7113 10421 7147 10455
rect 8033 10421 8067 10455
rect 11713 10421 11747 10455
rect 15117 10421 15151 10455
rect 6311 10217 6345 10251
rect 9781 10217 9815 10251
rect 12725 10217 12759 10251
rect 13293 10217 13327 10251
rect 13461 10217 13495 10251
rect 5441 10149 5475 10183
rect 5641 10149 5675 10183
rect 6101 10149 6135 10183
rect 7481 10149 7515 10183
rect 9229 10149 9263 10183
rect 12449 10149 12483 10183
rect 13093 10149 13127 10183
rect 6745 10081 6779 10115
rect 7113 10081 7147 10115
rect 9689 10081 9723 10115
rect 10333 10081 10367 10115
rect 10517 10081 10551 10115
rect 10977 10081 11011 10115
rect 12633 10081 12667 10115
rect 12817 10081 12851 10115
rect 13553 10081 13587 10115
rect 14381 10081 14415 10115
rect 6561 10013 6595 10047
rect 9965 10013 9999 10047
rect 14105 10013 14139 10047
rect 7297 9945 7331 9979
rect 13001 9945 13035 9979
rect 5273 9877 5307 9911
rect 5457 9877 5491 9911
rect 6285 9877 6319 9911
rect 6469 9877 6503 9911
rect 6929 9877 6963 9911
rect 9321 9877 9355 9911
rect 10149 9877 10183 9911
rect 11069 9877 11103 9911
rect 13277 9877 13311 9911
rect 13737 9877 13771 9911
rect 15669 9877 15703 9911
rect 5825 9673 5859 9707
rect 8677 9673 8711 9707
rect 10425 9673 10459 9707
rect 10609 9673 10643 9707
rect 11897 9673 11931 9707
rect 6653 9605 6687 9639
rect 9965 9605 9999 9639
rect 10977 9605 11011 9639
rect 12817 9605 12851 9639
rect 12909 9605 12943 9639
rect 4445 9537 4479 9571
rect 8953 9537 8987 9571
rect 9045 9537 9079 9571
rect 9413 9537 9447 9571
rect 10149 9537 10183 9571
rect 12173 9537 12207 9571
rect 12633 9537 12667 9571
rect 6009 9469 6043 9503
rect 8033 9469 8067 9503
rect 9321 9469 9355 9503
rect 10057 9469 10091 9503
rect 10701 9469 10735 9503
rect 12541 9469 12575 9503
rect 13139 9469 13173 9503
rect 13369 9469 13403 9503
rect 13737 9469 13771 9503
rect 4712 9401 4746 9435
rect 6561 9401 6595 9435
rect 7766 9401 7800 9435
rect 8493 9401 8527 9435
rect 8698 9401 8732 9435
rect 9689 9401 9723 9435
rect 10241 9401 10275 9435
rect 10977 9401 11011 9435
rect 11713 9401 11747 9435
rect 12265 9401 12299 9435
rect 13982 9401 14016 9435
rect 8861 9333 8895 9367
rect 9229 9333 9263 9367
rect 9597 9333 9631 9367
rect 9781 9333 9815 9367
rect 10441 9333 10475 9367
rect 10793 9333 10827 9367
rect 11913 9333 11947 9367
rect 12081 9333 12115 9367
rect 13277 9333 13311 9367
rect 15117 9333 15151 9367
rect 4997 9129 5031 9163
rect 5917 9129 5951 9163
rect 7389 9129 7423 9163
rect 9965 9129 9999 9163
rect 12173 9129 12207 9163
rect 13461 9129 13495 9163
rect 13737 9129 13771 9163
rect 6469 9061 6503 9095
rect 6561 9061 6595 9095
rect 10149 9061 10183 9095
rect 14096 9061 14130 9095
rect 5181 8993 5215 9027
rect 6193 8993 6227 9027
rect 6653 8993 6687 9027
rect 6837 8993 6871 9027
rect 7205 8993 7239 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 9873 8993 9907 9027
rect 10333 8993 10367 9027
rect 12449 8993 12483 9027
rect 12725 8993 12759 9027
rect 13093 8993 13127 9027
rect 13277 8993 13311 9027
rect 13553 8993 13587 9027
rect 6101 8925 6135 8959
rect 6929 8925 6963 8959
rect 7021 8925 7055 8959
rect 12357 8925 12391 8959
rect 12817 8925 12851 8959
rect 13001 8925 13035 8959
rect 13185 8925 13219 8959
rect 13829 8925 13863 8959
rect 9229 8789 9263 8823
rect 15209 8789 15243 8823
rect 5825 8585 5859 8619
rect 10333 8585 10367 8619
rect 12541 8585 12575 8619
rect 12357 8517 12391 8551
rect 6009 8381 6043 8415
rect 6193 8381 6227 8415
rect 6285 8381 6319 8415
rect 6561 8381 6595 8415
rect 6745 8381 6779 8415
rect 6837 8381 6871 8415
rect 8769 8381 8803 8415
rect 8953 8381 8987 8415
rect 9229 8381 9263 8415
rect 10885 8381 10919 8415
rect 11069 8381 11103 8415
rect 11253 8381 11287 8415
rect 12725 8313 12759 8347
rect 6377 8245 6411 8279
rect 9413 8245 9447 8279
rect 11161 8245 11195 8279
rect 12525 8245 12559 8279
rect 9965 8041 9999 8075
rect 10977 8041 11011 8075
rect 8401 7973 8435 8007
rect 9781 7973 9815 8007
rect 10333 7973 10367 8007
rect 12541 7973 12575 8007
rect 6009 7905 6043 7939
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 6561 7905 6595 7939
rect 7573 7905 7607 7939
rect 8309 7905 8343 7939
rect 8769 7905 8803 7939
rect 9045 7905 9079 7939
rect 9137 7905 9171 7939
rect 9321 7905 9355 7939
rect 9413 7905 9447 7939
rect 9597 7905 9631 7939
rect 11345 7905 11379 7939
rect 11989 7905 12023 7939
rect 12173 7905 12207 7939
rect 12449 7905 12483 7939
rect 12725 7905 12759 7939
rect 12909 7905 12943 7939
rect 13093 7905 13127 7939
rect 7113 7837 7147 7871
rect 7481 7837 7515 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8953 7837 8987 7871
rect 10425 7837 10459 7871
rect 10609 7837 10643 7871
rect 11437 7837 11471 7871
rect 11529 7837 11563 7871
rect 7297 7769 7331 7803
rect 13001 7769 13035 7803
rect 5825 7701 5859 7735
rect 7941 7701 7975 7735
rect 8125 7701 8159 7735
rect 8585 7701 8619 7735
rect 12357 7701 12391 7735
rect 12725 7701 12759 7735
rect 7113 7497 7147 7531
rect 10977 7497 11011 7531
rect 6285 7361 6319 7395
rect 6561 7361 6595 7395
rect 8401 7361 8435 7395
rect 8677 7361 8711 7395
rect 12357 7361 12391 7395
rect 6653 7293 6687 7327
rect 6929 7293 6963 7327
rect 7297 7293 7331 7327
rect 12090 7293 12124 7327
rect 12449 7293 12483 7327
rect 12633 7293 12667 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 13001 7293 13035 7327
rect 4905 7225 4939 7259
rect 6745 7157 6779 7191
rect 7941 7157 7975 7191
rect 9781 7157 9815 7191
rect 13185 7157 13219 7191
rect 8861 6953 8895 6987
rect 12357 6953 12391 6987
rect 8217 6885 8251 6919
rect 8417 6885 8451 6919
rect 13470 6885 13504 6919
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 8677 6817 8711 6851
rect 8953 6817 8987 6851
rect 9413 6817 9447 6851
rect 13737 6817 13771 6851
rect 9137 6749 9171 6783
rect 8677 6681 8711 6715
rect 6561 6613 6595 6647
rect 8401 6613 8435 6647
rect 8585 6613 8619 6647
rect 10701 6613 10735 6647
rect 9321 6273 9355 6307
rect 9597 6273 9631 6307
rect 10977 6137 11011 6171
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 9490 18884 9496 18896
rect 8956 18856 9496 18884
rect 842 18776 848 18828
rect 900 18816 906 18828
rect 937 18819 995 18825
rect 937 18816 949 18819
rect 900 18788 949 18816
rect 900 18776 906 18788
rect 937 18785 949 18788
rect 983 18785 995 18819
rect 937 18779 995 18785
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 2593 18819 2651 18825
rect 2593 18816 2605 18819
rect 2556 18788 2605 18816
rect 2556 18776 2562 18788
rect 2593 18785 2605 18788
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4212 18788 4261 18816
rect 4212 18776 4218 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5868 18788 5917 18816
rect 5868 18776 5874 18788
rect 5905 18785 5917 18788
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 8956 18825 8984 18856
rect 9490 18844 9496 18856
rect 9548 18844 9554 18896
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7524 18788 7573 18816
rect 7524 18776 7530 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 8941 18819 8999 18825
rect 8941 18785 8953 18819
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9585 18819 9643 18825
rect 9585 18816 9597 18819
rect 9180 18788 9597 18816
rect 9180 18776 9186 18788
rect 9585 18785 9597 18788
rect 9631 18785 9643 18819
rect 9585 18779 9643 18785
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 10965 18819 11023 18825
rect 10965 18816 10977 18819
rect 10836 18788 10977 18816
rect 10836 18776 10842 18788
rect 10965 18785 10977 18788
rect 11011 18785 11023 18819
rect 10965 18779 11023 18785
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12492 18788 12725 18816
rect 12492 18776 12498 18788
rect 12713 18785 12725 18788
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14148 18788 14381 18816
rect 14148 18776 14154 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15804 18788 16313 18816
rect 15804 18776 15810 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17460 18788 17693 18816
rect 17460 18776 17466 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 1213 18751 1271 18757
rect 1213 18717 1225 18751
rect 1259 18748 1271 18751
rect 6914 18748 6920 18760
rect 1259 18720 6920 18748
rect 1259 18717 1271 18720
rect 1213 18711 1271 18717
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 8849 18751 8907 18757
rect 8849 18717 8861 18751
rect 8895 18717 8907 18751
rect 8849 18711 8907 18717
rect 2777 18683 2835 18689
rect 2777 18649 2789 18683
rect 2823 18680 2835 18683
rect 6270 18680 6276 18692
rect 2823 18652 6276 18680
rect 2823 18649 2835 18652
rect 2777 18643 2835 18649
rect 6270 18640 6276 18652
rect 6328 18640 6334 18692
rect 8864 18680 8892 18711
rect 9306 18708 9312 18760
rect 9364 18708 9370 18760
rect 8864 18652 9444 18680
rect 9416 18624 9444 18652
rect 13170 18640 13176 18692
rect 13228 18680 13234 18692
rect 16117 18683 16175 18689
rect 16117 18680 16129 18683
rect 13228 18652 16129 18680
rect 13228 18640 13234 18652
rect 16117 18649 16129 18652
rect 16163 18649 16175 18683
rect 16117 18643 16175 18649
rect 4433 18615 4491 18621
rect 4433 18581 4445 18615
rect 4479 18612 4491 18615
rect 5902 18612 5908 18624
rect 4479 18584 5908 18612
rect 4479 18581 4491 18584
rect 4433 18575 4491 18581
rect 5902 18572 5908 18584
rect 5960 18572 5966 18624
rect 6089 18615 6147 18621
rect 6089 18581 6101 18615
rect 6135 18612 6147 18615
rect 6638 18612 6644 18624
rect 6135 18584 6644 18612
rect 6135 18581 6147 18584
rect 6089 18575 6147 18581
rect 6638 18572 6644 18584
rect 6696 18572 6702 18624
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 8570 18612 8576 18624
rect 7791 18584 8576 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8662 18572 8668 18624
rect 8720 18572 8726 18624
rect 9398 18572 9404 18624
rect 9456 18572 9462 18624
rect 10870 18572 10876 18624
rect 10928 18612 10934 18624
rect 11149 18615 11207 18621
rect 11149 18612 11161 18615
rect 10928 18584 11161 18612
rect 10928 18572 10934 18584
rect 11149 18581 11161 18584
rect 11195 18581 11207 18615
rect 11149 18575 11207 18581
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 14182 18572 14188 18624
rect 14240 18572 14246 18624
rect 17494 18572 17500 18624
rect 17552 18572 17558 18624
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 7101 18411 7159 18417
rect 7101 18377 7113 18411
rect 7147 18408 7159 18411
rect 9490 18408 9496 18420
rect 7147 18380 9496 18408
rect 7147 18377 7159 18380
rect 7101 18371 7159 18377
rect 9490 18368 9496 18380
rect 9548 18368 9554 18420
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18309 6883 18343
rect 6825 18303 6883 18309
rect 9769 18343 9827 18349
rect 9769 18309 9781 18343
rect 9815 18309 9827 18343
rect 9769 18303 9827 18309
rect 6840 18272 6868 18303
rect 6840 18244 7328 18272
rect 5442 18164 5448 18216
rect 5500 18164 5506 18216
rect 6914 18164 6920 18216
rect 6972 18164 6978 18216
rect 7300 18213 7328 18244
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 8386 18164 8392 18216
rect 8444 18164 8450 18216
rect 8662 18213 8668 18216
rect 8656 18204 8668 18213
rect 8623 18176 8668 18204
rect 8656 18167 8668 18176
rect 8662 18164 8668 18167
rect 8720 18164 8726 18216
rect 9784 18204 9812 18303
rect 13004 18244 13308 18272
rect 13004 18216 13032 18244
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9784 18176 9873 18204
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 9861 18167 9919 18173
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 12986 18204 12992 18216
rect 11112 18176 12992 18204
rect 11112 18164 11118 18176
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 13078 18164 13084 18216
rect 13136 18164 13142 18216
rect 13170 18164 13176 18216
rect 13228 18164 13234 18216
rect 13280 18204 13308 18244
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 13280 18176 14933 18204
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 15105 18207 15163 18213
rect 15105 18204 15117 18207
rect 14967 18176 15117 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 15105 18173 15117 18176
rect 15151 18173 15163 18207
rect 15105 18167 15163 18173
rect 17129 18207 17187 18213
rect 17129 18173 17141 18207
rect 17175 18204 17187 18207
rect 17494 18204 17500 18216
rect 17175 18176 17500 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 5712 18139 5770 18145
rect 5712 18105 5724 18139
rect 5758 18136 5770 18139
rect 5994 18136 6000 18148
rect 5758 18108 6000 18136
rect 5758 18105 5770 18108
rect 5712 18099 5770 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 11324 18139 11382 18145
rect 11324 18105 11336 18139
rect 11370 18136 11382 18139
rect 12342 18136 12348 18148
rect 11370 18108 12348 18136
rect 11370 18105 11382 18108
rect 11324 18099 11382 18105
rect 12342 18096 12348 18108
rect 12400 18096 12406 18148
rect 13357 18139 13415 18145
rect 13357 18105 13369 18139
rect 13403 18136 13415 18139
rect 14654 18139 14712 18145
rect 14654 18136 14666 18139
rect 13403 18108 14666 18136
rect 13403 18105 13415 18108
rect 13357 18099 13415 18105
rect 14654 18105 14666 18108
rect 14700 18105 14712 18139
rect 14654 18099 14712 18105
rect 15378 18096 15384 18148
rect 15436 18096 15442 18148
rect 17037 18139 17095 18145
rect 17037 18136 17049 18139
rect 16606 18108 17049 18136
rect 17037 18105 17049 18108
rect 17083 18105 17095 18139
rect 17037 18099 17095 18105
rect 7374 18028 7380 18080
rect 7432 18028 7438 18080
rect 9214 18028 9220 18080
rect 9272 18068 9278 18080
rect 9953 18071 10011 18077
rect 9953 18068 9965 18071
rect 9272 18040 9965 18068
rect 9272 18028 9278 18040
rect 9953 18037 9965 18040
rect 9999 18037 10011 18071
rect 9953 18031 10011 18037
rect 12434 18028 12440 18080
rect 12492 18028 12498 18080
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 13541 18071 13599 18077
rect 13541 18037 13553 18071
rect 13587 18068 13599 18071
rect 13722 18068 13728 18080
rect 13587 18040 13728 18068
rect 13587 18037 13599 18040
rect 13541 18031 13599 18037
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 16666 18028 16672 18080
rect 16724 18068 16730 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 16724 18040 16865 18068
rect 16724 18028 16730 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 5994 17824 6000 17876
rect 6052 17824 6058 17876
rect 6641 17867 6699 17873
rect 6641 17833 6653 17867
rect 6687 17864 6699 17867
rect 6733 17867 6791 17873
rect 6733 17864 6745 17867
rect 6687 17836 6745 17864
rect 6687 17833 6699 17836
rect 6641 17827 6699 17833
rect 6733 17833 6745 17836
rect 6779 17833 6791 17867
rect 6733 17827 6791 17833
rect 8849 17867 8907 17873
rect 8849 17833 8861 17867
rect 8895 17864 8907 17867
rect 9306 17864 9312 17876
rect 8895 17836 9312 17864
rect 8895 17833 8907 17836
rect 8849 17827 8907 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 12342 17824 12348 17876
rect 12400 17824 12406 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 12989 17867 13047 17873
rect 12989 17864 13001 17867
rect 12768 17836 13001 17864
rect 12768 17824 12774 17836
rect 12989 17833 13001 17836
rect 13035 17833 13047 17867
rect 12989 17827 13047 17833
rect 15378 17824 15384 17876
rect 15436 17864 15442 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 15436 17836 15485 17864
rect 15436 17824 15442 17836
rect 15473 17833 15485 17836
rect 15519 17833 15531 17867
rect 15473 17827 15531 17833
rect 8386 17796 8392 17808
rect 7392 17768 8392 17796
rect 5902 17688 5908 17740
rect 5960 17728 5966 17740
rect 6273 17731 6331 17737
rect 6273 17728 6285 17731
rect 5960 17700 6285 17728
rect 5960 17688 5966 17700
rect 6273 17697 6285 17700
rect 6319 17697 6331 17731
rect 6273 17691 6331 17697
rect 6914 17688 6920 17740
rect 6972 17688 6978 17740
rect 7101 17731 7159 17737
rect 7101 17697 7113 17731
rect 7147 17728 7159 17731
rect 7282 17728 7288 17740
rect 7147 17700 7288 17728
rect 7147 17697 7159 17700
rect 7101 17691 7159 17697
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 6181 17663 6239 17669
rect 6181 17629 6193 17663
rect 6227 17660 6239 17663
rect 6546 17660 6552 17672
rect 6227 17632 6552 17660
rect 6227 17629 6239 17632
rect 6181 17623 6239 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 7392 17669 7420 17768
rect 8386 17756 8392 17768
rect 8444 17796 8450 17808
rect 8444 17768 9444 17796
rect 8444 17756 8450 17768
rect 7644 17731 7702 17737
rect 7644 17697 7656 17731
rect 7690 17728 7702 17731
rect 9030 17728 9036 17740
rect 7690 17700 9036 17728
rect 7690 17697 7702 17700
rect 7644 17691 7702 17697
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 9416 17737 9444 17768
rect 9490 17756 9496 17808
rect 9548 17796 9554 17808
rect 9548 17768 11284 17796
rect 9548 17756 9554 17768
rect 11256 17737 11284 17768
rect 12084 17768 13124 17796
rect 12084 17737 12112 17768
rect 13096 17740 13124 17768
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 13228 17768 13676 17796
rect 13228 17756 13234 17768
rect 9217 17731 9275 17737
rect 9217 17697 9229 17731
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 9401 17731 9459 17737
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9668 17731 9726 17737
rect 9668 17697 9680 17731
rect 9714 17728 9726 17731
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 9714 17700 10977 17728
rect 9714 17697 9726 17700
rect 9668 17691 9726 17697
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 11241 17731 11299 17737
rect 11241 17697 11253 17731
rect 11287 17728 11299 17731
rect 12069 17731 12127 17737
rect 12069 17728 12081 17731
rect 11287 17700 12081 17728
rect 11287 17697 11299 17700
rect 11241 17691 11299 17697
rect 12069 17697 12081 17700
rect 12115 17697 12127 17731
rect 12069 17691 12127 17697
rect 7377 17663 7435 17669
rect 7377 17629 7389 17663
rect 7423 17629 7435 17663
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 7377 17623 7435 17629
rect 8404 17632 9137 17660
rect 5442 17552 5448 17604
rect 5500 17592 5506 17604
rect 7392 17592 7420 17623
rect 5500 17564 7420 17592
rect 5500 17552 5506 17564
rect 7101 17527 7159 17533
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7374 17524 7380 17536
rect 7147 17496 7380 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8404 17524 8432 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 8478 17552 8484 17604
rect 8536 17592 8542 17604
rect 9232 17592 9260 17691
rect 12434 17688 12440 17740
rect 12492 17688 12498 17740
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13265 17731 13323 17737
rect 13265 17728 13277 17731
rect 13136 17700 13277 17728
rect 13136 17688 13142 17700
rect 13265 17697 13277 17700
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 13354 17688 13360 17740
rect 13412 17688 13418 17740
rect 13648 17737 13676 17768
rect 13633 17731 13691 17737
rect 13633 17697 13645 17731
rect 13679 17697 13691 17731
rect 13633 17691 13691 17697
rect 13722 17688 13728 17740
rect 13780 17688 13786 17740
rect 10870 17620 10876 17672
rect 10928 17660 10934 17672
rect 11149 17663 11207 17669
rect 11149 17660 11161 17663
rect 10928 17632 11161 17660
rect 10928 17620 10934 17632
rect 11149 17629 11161 17632
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 9306 17592 9312 17604
rect 8536 17564 9312 17592
rect 8536 17552 8542 17564
rect 9306 17552 9312 17564
rect 9364 17552 9370 17604
rect 10502 17552 10508 17604
rect 10560 17592 10566 17604
rect 11624 17592 11652 17623
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17660 12219 17663
rect 12526 17660 12532 17672
rect 12207 17632 12532 17660
rect 12207 17629 12219 17632
rect 12161 17623 12219 17629
rect 12526 17620 12532 17632
rect 12584 17620 12590 17672
rect 10560 17564 11652 17592
rect 13372 17564 13860 17592
rect 10560 17552 10566 17564
rect 8168 17496 8432 17524
rect 8168 17484 8174 17496
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8720 17496 8769 17524
rect 8720 17484 8726 17496
rect 8757 17493 8769 17496
rect 8803 17493 8815 17527
rect 8757 17487 8815 17493
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 9582 17524 9588 17536
rect 9272 17496 9588 17524
rect 9272 17484 9278 17496
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 10781 17527 10839 17533
rect 10781 17493 10793 17527
rect 10827 17524 10839 17527
rect 11606 17524 11612 17536
rect 10827 17496 11612 17524
rect 10827 17493 10839 17496
rect 10781 17487 10839 17493
rect 11606 17484 11612 17496
rect 11664 17484 11670 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12618 17524 12624 17536
rect 12575 17496 12624 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 13372 17533 13400 17564
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 13541 17527 13599 17533
rect 13541 17493 13553 17527
rect 13587 17524 13599 17527
rect 13630 17524 13636 17536
rect 13587 17496 13636 17524
rect 13587 17493 13599 17496
rect 13541 17487 13599 17493
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 13832 17533 13860 17564
rect 13817 17527 13875 17533
rect 13817 17493 13829 17527
rect 13863 17524 13875 17527
rect 13998 17524 14004 17536
rect 13863 17496 14004 17524
rect 13863 17493 13875 17496
rect 13817 17487 13875 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 7190 17280 7196 17332
rect 7248 17280 7254 17332
rect 8021 17323 8079 17329
rect 8021 17289 8033 17323
rect 8067 17320 8079 17323
rect 8938 17320 8944 17332
rect 8067 17292 8944 17320
rect 8067 17289 8079 17292
rect 8021 17283 8079 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9030 17280 9036 17332
rect 9088 17280 9094 17332
rect 10318 17280 10324 17332
rect 10376 17280 10382 17332
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 10965 17323 11023 17329
rect 10965 17289 10977 17323
rect 11011 17289 11023 17323
rect 10965 17283 11023 17289
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 11698 17320 11704 17332
rect 11287 17292 11704 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 10980 17252 11008 17283
rect 11698 17280 11704 17292
rect 11756 17280 11762 17332
rect 16666 17320 16672 17332
rect 12728 17292 16672 17320
rect 12618 17252 12624 17264
rect 8128 17224 10272 17252
rect 10980 17224 12624 17252
rect 8128 17196 8156 17224
rect 6457 17187 6515 17193
rect 6457 17153 6469 17187
rect 6503 17184 6515 17187
rect 6638 17184 6644 17196
rect 6503 17156 6644 17184
rect 6503 17153 6515 17156
rect 6457 17147 6515 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7208 17156 7941 17184
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4801 17119 4859 17125
rect 4801 17116 4813 17119
rect 4212 17088 4813 17116
rect 4212 17076 4218 17088
rect 4801 17085 4813 17088
rect 4847 17116 4859 17119
rect 5442 17116 5448 17128
rect 4847 17088 5448 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 6546 17076 6552 17128
rect 6604 17076 6610 17128
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7208 17125 7236 17156
rect 7929 17153 7941 17156
rect 7975 17184 7987 17187
rect 8110 17184 8116 17196
rect 7975 17156 8116 17184
rect 7975 17153 7987 17156
rect 7929 17147 7987 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8849 17187 8907 17193
rect 8849 17184 8861 17187
rect 8628 17156 8861 17184
rect 8628 17144 8634 17156
rect 8849 17153 8861 17156
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 7193 17119 7251 17125
rect 7193 17116 7205 17119
rect 6972 17088 7205 17116
rect 6972 17076 6978 17088
rect 7193 17085 7205 17088
rect 7239 17085 7251 17119
rect 7193 17079 7251 17085
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7377 17119 7435 17125
rect 7377 17116 7389 17119
rect 7340 17088 7389 17116
rect 7340 17076 7346 17088
rect 7377 17085 7389 17088
rect 7423 17116 7435 17119
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7423 17088 7849 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 7837 17085 7849 17088
rect 7883 17116 7895 17119
rect 8018 17116 8024 17128
rect 7883 17088 8024 17116
rect 7883 17085 7895 17088
rect 7837 17079 7895 17085
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17085 8815 17119
rect 8864 17116 8892 17147
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 10244 17193 10272 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 10229 17187 10287 17193
rect 9364 17156 10180 17184
rect 9364 17144 9370 17156
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 8864 17088 9137 17116
rect 8757 17079 8815 17085
rect 9125 17085 9137 17088
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 5068 17051 5126 17057
rect 5068 17017 5080 17051
rect 5114 17048 5126 17051
rect 6273 17051 6331 17057
rect 6273 17048 6285 17051
rect 5114 17020 6285 17048
rect 5114 17017 5126 17020
rect 5068 17011 5126 17017
rect 6273 17017 6285 17020
rect 6319 17017 6331 17051
rect 6564 17048 6592 17076
rect 8772 17048 8800 17079
rect 9490 17076 9496 17128
rect 9548 17076 9554 17128
rect 10152 17125 10180 17156
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10275 17156 10977 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 12526 17184 12532 17196
rect 10965 17147 11023 17153
rect 11532 17156 12532 17184
rect 10137 17119 10195 17125
rect 10137 17085 10149 17119
rect 10183 17116 10195 17119
rect 10873 17119 10931 17125
rect 10873 17116 10885 17119
rect 10183 17088 10885 17116
rect 10183 17085 10195 17088
rect 10137 17079 10195 17085
rect 10873 17085 10885 17088
rect 10919 17116 10931 17119
rect 11422 17116 11428 17128
rect 10919 17088 11428 17116
rect 10919 17085 10931 17088
rect 10873 17079 10931 17085
rect 11422 17076 11428 17088
rect 11480 17076 11486 17128
rect 11532 17125 11560 17156
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11606 17076 11612 17128
rect 11664 17076 11670 17128
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 12728 17116 12756 17292
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13538 17184 13544 17196
rect 13044 17156 13544 17184
rect 13044 17144 13050 17156
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 12216 17088 12756 17116
rect 12216 17076 12222 17088
rect 13078 17076 13084 17128
rect 13136 17076 13142 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 14182 17116 14188 17128
rect 13228 17088 14188 17116
rect 13228 17076 13234 17088
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 9508 17048 9536 17076
rect 6564 17020 9536 17048
rect 6273 17011 6331 17017
rect 10318 17008 10324 17060
rect 10376 17048 10382 17060
rect 10778 17048 10784 17060
rect 10376 17020 10784 17048
rect 10376 17008 10382 17020
rect 10778 17008 10784 17020
rect 10836 17048 10842 17060
rect 11701 17051 11759 17057
rect 11701 17048 11713 17051
rect 10836 17020 11713 17048
rect 10836 17008 10842 17020
rect 11701 17017 11713 17020
rect 11747 17017 11759 17051
rect 11701 17011 11759 17017
rect 13357 17051 13415 17057
rect 13357 17017 13369 17051
rect 13403 17048 13415 17051
rect 13786 17051 13844 17057
rect 13786 17048 13798 17051
rect 13403 17020 13798 17048
rect 13403 17017 13415 17020
rect 13357 17011 13415 17017
rect 13786 17017 13798 17020
rect 13832 17017 13844 17051
rect 13786 17011 13844 17017
rect 6181 16983 6239 16989
rect 6181 16949 6193 16983
rect 6227 16980 6239 16983
rect 6362 16980 6368 16992
rect 6227 16952 6368 16980
rect 6227 16949 6239 16952
rect 6181 16943 6239 16949
rect 6362 16940 6368 16952
rect 6420 16940 6426 16992
rect 6917 16983 6975 16989
rect 6917 16949 6929 16983
rect 6963 16980 6975 16983
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 6963 16952 7021 16980
rect 6963 16949 6975 16952
rect 6917 16943 6975 16949
rect 7009 16949 7021 16952
rect 7055 16949 7067 16983
rect 7009 16943 7067 16949
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8389 16983 8447 16989
rect 8389 16980 8401 16983
rect 8251 16952 8401 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8389 16949 8401 16952
rect 8435 16949 8447 16983
rect 8389 16943 8447 16949
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9490 16980 9496 16992
rect 9263 16952 9496 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 11330 16940 11336 16992
rect 11388 16980 11394 16992
rect 11425 16983 11483 16989
rect 11425 16980 11437 16983
rect 11388 16952 11437 16980
rect 11388 16940 11394 16952
rect 11425 16949 11437 16952
rect 11471 16949 11483 16983
rect 11425 16943 11483 16949
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 12342 16980 12348 16992
rect 11572 16952 12348 16980
rect 11572 16940 11578 16952
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 12713 16983 12771 16989
rect 12713 16949 12725 16983
rect 12759 16980 12771 16983
rect 12894 16980 12900 16992
rect 12759 16952 12900 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 13906 16940 13912 16992
rect 13964 16980 13970 16992
rect 14921 16983 14979 16989
rect 14921 16980 14933 16983
rect 13964 16952 14933 16980
rect 13964 16940 13970 16952
rect 14921 16949 14933 16952
rect 14967 16949 14979 16983
rect 14921 16943 14979 16949
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 6696 16748 7972 16776
rect 6696 16736 6702 16748
rect 6457 16711 6515 16717
rect 6457 16677 6469 16711
rect 6503 16708 6515 16711
rect 6503 16680 7052 16708
rect 6503 16677 6515 16680
rect 6457 16671 6515 16677
rect 6362 16600 6368 16652
rect 6420 16600 6426 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 6656 16504 6684 16603
rect 6914 16600 6920 16652
rect 6972 16600 6978 16652
rect 7024 16649 7052 16680
rect 7009 16643 7067 16649
rect 7009 16609 7021 16643
rect 7055 16640 7067 16643
rect 7190 16640 7196 16652
rect 7055 16612 7196 16640
rect 7055 16609 7067 16612
rect 7009 16603 7067 16609
rect 7190 16600 7196 16612
rect 7248 16640 7254 16652
rect 7834 16640 7840 16652
rect 7248 16612 7840 16640
rect 7248 16600 7254 16612
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 7944 16640 7972 16748
rect 8938 16736 8944 16788
rect 8996 16776 9002 16788
rect 9309 16779 9367 16785
rect 9309 16776 9321 16779
rect 8996 16748 9321 16776
rect 8996 16736 9002 16748
rect 9309 16745 9321 16748
rect 9355 16745 9367 16779
rect 9309 16739 9367 16745
rect 12894 16736 12900 16788
rect 12952 16736 12958 16788
rect 8018 16668 8024 16720
rect 8076 16708 8082 16720
rect 12158 16708 12164 16720
rect 8076 16680 12164 16708
rect 8076 16668 8082 16680
rect 12158 16668 12164 16680
rect 12216 16668 12222 16720
rect 7944 16612 8616 16640
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 7374 16572 7380 16584
rect 6779 16544 7380 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 7374 16532 7380 16544
rect 7432 16532 7438 16584
rect 8588 16572 8616 16612
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 9217 16643 9275 16649
rect 9217 16640 9229 16643
rect 8720 16612 9229 16640
rect 8720 16600 8726 16612
rect 9217 16609 9229 16612
rect 9263 16609 9275 16643
rect 10594 16640 10600 16652
rect 9217 16603 9275 16609
rect 9324 16612 10600 16640
rect 9324 16572 9352 16612
rect 10594 16600 10600 16612
rect 10652 16600 10658 16652
rect 12342 16600 12348 16652
rect 12400 16640 12406 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12400 16612 13277 16640
rect 12400 16600 12406 16612
rect 13265 16609 13277 16612
rect 13311 16640 13323 16643
rect 13354 16640 13360 16652
rect 13311 16612 13360 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13906 16600 13912 16652
rect 13964 16600 13970 16652
rect 8588 16544 9352 16572
rect 13078 16532 13084 16584
rect 13136 16572 13142 16584
rect 13173 16575 13231 16581
rect 13173 16572 13185 16575
rect 13136 16544 13185 16572
rect 13136 16532 13142 16544
rect 13173 16541 13185 16544
rect 13219 16541 13231 16575
rect 13173 16535 13231 16541
rect 7006 16504 7012 16516
rect 6656 16476 7012 16504
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 7190 16396 7196 16448
rect 7248 16396 7254 16448
rect 8846 16396 8852 16448
rect 8904 16396 8910 16448
rect 9125 16439 9183 16445
rect 9125 16405 9137 16439
rect 9171 16436 9183 16439
rect 9214 16436 9220 16448
rect 9171 16408 9220 16436
rect 9171 16405 9183 16408
rect 9125 16399 9183 16405
rect 9214 16396 9220 16408
rect 9272 16396 9278 16448
rect 13265 16439 13323 16445
rect 13265 16405 13277 16439
rect 13311 16436 13323 16439
rect 13814 16436 13820 16448
rect 13311 16408 13820 16436
rect 13311 16405 13323 16408
rect 13265 16399 13323 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 6914 16232 6920 16244
rect 6840 16204 6920 16232
rect 6457 16167 6515 16173
rect 6457 16133 6469 16167
rect 6503 16164 6515 16167
rect 6638 16164 6644 16176
rect 6503 16136 6644 16164
rect 6503 16133 6515 16136
rect 6457 16127 6515 16133
rect 6638 16124 6644 16136
rect 6696 16124 6702 16176
rect 6181 16031 6239 16037
rect 6181 15997 6193 16031
rect 6227 15997 6239 16031
rect 6181 15991 6239 15997
rect 6196 15960 6224 15991
rect 6270 15988 6276 16040
rect 6328 16028 6334 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6328 16000 6653 16028
rect 6328 15988 6334 16000
rect 6641 15997 6653 16000
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6730 15988 6736 16040
rect 6788 16037 6794 16040
rect 6840 16037 6868 16204
rect 6914 16192 6920 16204
rect 6972 16232 6978 16244
rect 7926 16232 7932 16244
rect 6972 16204 7932 16232
rect 6972 16192 6978 16204
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 10318 16232 10324 16244
rect 9416 16204 10324 16232
rect 9416 16173 9444 16204
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 7285 16167 7343 16173
rect 7285 16133 7297 16167
rect 7331 16133 7343 16167
rect 7285 16127 7343 16133
rect 9401 16167 9459 16173
rect 9401 16133 9413 16167
rect 9447 16133 9459 16167
rect 11146 16164 11152 16176
rect 9401 16127 9459 16133
rect 9600 16136 11152 16164
rect 7300 16096 7328 16127
rect 9306 16096 9312 16108
rect 7300 16068 8800 16096
rect 6788 16031 6868 16037
rect 6788 15997 6801 16031
rect 6835 16000 6868 16031
rect 6835 15997 6847 16000
rect 6788 15991 6847 15997
rect 6788 15988 6794 15991
rect 7006 15988 7012 16040
rect 7064 15988 7070 16040
rect 7147 16031 7205 16037
rect 7147 15997 7159 16031
rect 7193 16028 7205 16031
rect 7374 16028 7380 16040
rect 7193 16000 7380 16028
rect 7193 15997 7205 16000
rect 7147 15991 7205 15997
rect 7374 15988 7380 16000
rect 7432 16028 7438 16040
rect 7561 16031 7619 16037
rect 7561 16028 7573 16031
rect 7432 16000 7573 16028
rect 7432 15988 7438 16000
rect 7561 15997 7573 16000
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 16028 7803 16031
rect 7834 16028 7840 16040
rect 7791 16000 7840 16028
rect 7791 15997 7803 16000
rect 7745 15991 7803 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8772 16037 8800 16068
rect 8864 16068 9312 16096
rect 8864 16037 8892 16068
rect 9306 16056 9312 16068
rect 9364 16056 9370 16108
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 15997 8907 16031
rect 8849 15991 8907 15997
rect 9214 15988 9220 16040
rect 9272 16028 9278 16040
rect 9493 16031 9551 16037
rect 9493 16028 9505 16031
rect 9272 16000 9505 16028
rect 9272 15988 9278 16000
rect 9493 15997 9505 16000
rect 9539 15997 9551 16031
rect 9493 15991 9551 15997
rect 6196 15932 6592 15960
rect 6089 15895 6147 15901
rect 6089 15861 6101 15895
rect 6135 15892 6147 15895
rect 6178 15892 6184 15904
rect 6135 15864 6184 15892
rect 6135 15861 6147 15864
rect 6089 15855 6147 15861
rect 6178 15852 6184 15864
rect 6236 15852 6242 15904
rect 6564 15892 6592 15932
rect 6914 15920 6920 15972
rect 6972 15920 6978 15972
rect 7024 15960 7052 15988
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 7024 15932 7665 15960
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 7653 15923 7711 15929
rect 9030 15920 9036 15972
rect 9088 15920 9094 15972
rect 9122 15920 9128 15972
rect 9180 15920 9186 15972
rect 9600 15960 9628 16136
rect 9692 16068 10824 16096
rect 9692 16037 9720 16068
rect 10796 16040 10824 16068
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 15997 9827 16031
rect 9769 15991 9827 15997
rect 9784 15960 9812 15991
rect 9858 15988 9864 16040
rect 9916 15988 9922 16040
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 16028 10103 16031
rect 10091 16000 10180 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 9600 15932 9812 15960
rect 7098 15892 7104 15904
rect 6564 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7374 15852 7380 15904
rect 7432 15852 7438 15904
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 10152 15892 10180 16000
rect 10778 15988 10784 16040
rect 10836 16028 10842 16040
rect 11072 16037 11100 16136
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 12618 16124 12624 16176
rect 12676 16124 12682 16176
rect 12636 16096 12664 16124
rect 12805 16099 12863 16105
rect 12805 16096 12817 16099
rect 11164 16068 12817 16096
rect 11164 16037 11192 16068
rect 12805 16065 12817 16068
rect 12851 16065 12863 16099
rect 12805 16059 12863 16065
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 13446 16096 13452 16108
rect 12943 16068 13452 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 13446 16056 13452 16068
rect 13504 16096 13510 16108
rect 13504 16068 13860 16096
rect 13504 16056 13510 16068
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10836 16000 10977 16028
rect 10836 15988 10842 16000
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11057 16031 11115 16037
rect 11057 15997 11069 16031
rect 11103 15997 11115 16031
rect 11057 15991 11115 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11333 16031 11391 16037
rect 11333 15997 11345 16031
rect 11379 16028 11391 16031
rect 12526 16028 12532 16040
rect 11379 16000 12532 16028
rect 11379 15997 11391 16000
rect 11333 15991 11391 15997
rect 12526 15988 12532 16000
rect 12584 16028 12590 16040
rect 12621 16031 12679 16037
rect 12621 16028 12633 16031
rect 12584 16000 12633 16028
rect 12584 15988 12590 16000
rect 12621 15997 12633 16000
rect 12667 15997 12679 16031
rect 12621 15991 12679 15997
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 15997 13047 16031
rect 12989 15991 13047 15997
rect 13173 16031 13231 16037
rect 13173 15997 13185 16031
rect 13219 16028 13231 16031
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 13219 16000 13553 16028
rect 13219 15997 13231 16000
rect 13173 15991 13231 15997
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 13004 15960 13032 15991
rect 13722 15988 13728 16040
rect 13780 15988 13786 16040
rect 13832 16037 13860 16068
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 13998 15988 14004 16040
rect 14056 15988 14062 16040
rect 14093 16031 14151 16037
rect 14093 15997 14105 16031
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 13740 15960 13768 15988
rect 13004 15932 13768 15960
rect 8628 15864 10180 15892
rect 8628 15852 8634 15864
rect 10226 15852 10232 15904
rect 10284 15852 10290 15904
rect 10502 15852 10508 15904
rect 10560 15892 10566 15904
rect 10781 15895 10839 15901
rect 10781 15892 10793 15895
rect 10560 15864 10793 15892
rect 10560 15852 10566 15864
rect 10781 15861 10793 15864
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 12434 15852 12440 15904
rect 12492 15852 12498 15904
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 14108 15892 14136 15991
rect 13044 15864 14136 15892
rect 13044 15852 13050 15864
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 6457 15691 6515 15697
rect 6457 15657 6469 15691
rect 6503 15688 6515 15691
rect 6914 15688 6920 15700
rect 6503 15660 6920 15688
rect 6503 15657 6515 15660
rect 6457 15651 6515 15657
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 7837 15691 7895 15697
rect 7837 15657 7849 15691
rect 7883 15688 7895 15691
rect 9030 15688 9036 15700
rect 7883 15660 9036 15688
rect 7883 15657 7895 15660
rect 7837 15651 7895 15657
rect 9030 15648 9036 15660
rect 9088 15648 9094 15700
rect 9122 15648 9128 15700
rect 9180 15688 9186 15700
rect 9180 15660 9628 15688
rect 9180 15648 9186 15660
rect 7282 15620 7288 15632
rect 6932 15592 7288 15620
rect 4516 15555 4574 15561
rect 4516 15521 4528 15555
rect 4562 15552 4574 15555
rect 5074 15552 5080 15564
rect 4562 15524 5080 15552
rect 4562 15521 4574 15524
rect 4516 15515 4574 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6932 15561 6960 15592
rect 7282 15580 7288 15592
rect 7340 15580 7346 15632
rect 7374 15580 7380 15632
rect 7432 15580 7438 15632
rect 8846 15580 8852 15632
rect 8904 15580 8910 15632
rect 6641 15555 6699 15561
rect 6641 15552 6653 15555
rect 6420 15524 6653 15552
rect 6420 15512 6426 15524
rect 6641 15521 6653 15524
rect 6687 15521 6699 15555
rect 6641 15515 6699 15521
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7006 15512 7012 15564
rect 7064 15552 7070 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 7064 15524 7113 15552
rect 7064 15512 7070 15524
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7101 15515 7159 15521
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 7116 15484 7144 15515
rect 8570 15512 8576 15564
rect 8628 15512 8634 15564
rect 8757 15555 8815 15561
rect 8757 15521 8769 15555
rect 8803 15521 8815 15555
rect 8757 15515 8815 15521
rect 7374 15484 7380 15496
rect 7116 15456 7380 15484
rect 4249 15447 4307 15453
rect 7374 15444 7380 15456
rect 7432 15444 7438 15496
rect 8772 15484 8800 15515
rect 8938 15512 8944 15564
rect 8996 15512 9002 15564
rect 9048 15552 9076 15648
rect 9600 15629 9628 15660
rect 13538 15648 13544 15700
rect 13596 15688 13602 15700
rect 14185 15691 14243 15697
rect 14185 15688 14197 15691
rect 13596 15660 14197 15688
rect 13596 15648 13602 15660
rect 14185 15657 14197 15660
rect 14231 15688 14243 15691
rect 14918 15688 14924 15700
rect 14231 15660 14924 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14918 15648 14924 15660
rect 14976 15648 14982 15700
rect 9585 15623 9643 15629
rect 9585 15589 9597 15623
rect 9631 15589 9643 15623
rect 12434 15620 12440 15632
rect 9585 15583 9643 15589
rect 10060 15592 10364 15620
rect 10060 15552 10088 15592
rect 10336 15561 10364 15592
rect 10428 15592 12440 15620
rect 10428 15561 10456 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 9048 15524 10088 15552
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10321 15555 10379 15561
rect 10321 15521 10333 15555
rect 10367 15521 10379 15555
rect 10321 15515 10379 15521
rect 10413 15555 10471 15561
rect 10413 15521 10425 15555
rect 10459 15521 10471 15555
rect 10413 15515 10471 15521
rect 9582 15484 9588 15496
rect 8772 15456 9588 15484
rect 9582 15444 9588 15456
rect 9640 15444 9646 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15484 10103 15487
rect 10152 15484 10180 15515
rect 10502 15512 10508 15564
rect 10560 15512 10566 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11221 15555 11279 15561
rect 11221 15552 11233 15555
rect 11112 15524 11233 15552
rect 11112 15512 11118 15524
rect 11221 15521 11233 15524
rect 11267 15521 11279 15555
rect 11221 15515 11279 15521
rect 12894 15512 12900 15564
rect 12952 15512 12958 15564
rect 10091 15456 10180 15484
rect 10091 15453 10103 15456
rect 10045 15447 10103 15453
rect 10962 15444 10968 15496
rect 11020 15444 11026 15496
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 7248 15388 7665 15416
rect 7248 15376 7254 15388
rect 7653 15385 7665 15388
rect 7699 15385 7711 15419
rect 7653 15379 7711 15385
rect 9953 15419 10011 15425
rect 9953 15385 9965 15419
rect 9999 15416 10011 15419
rect 10226 15416 10232 15428
rect 9999 15388 10232 15416
rect 9999 15385 10011 15388
rect 9953 15379 10011 15385
rect 10226 15376 10232 15388
rect 10284 15376 10290 15428
rect 5626 15308 5632 15360
rect 5684 15308 5690 15360
rect 9306 15308 9312 15360
rect 9364 15348 9370 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 9364 15320 10793 15348
rect 9364 15308 9370 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 12345 15351 12403 15357
rect 12345 15348 12357 15351
rect 11204 15320 12357 15348
rect 11204 15308 11210 15320
rect 12345 15317 12357 15320
rect 12391 15317 12403 15351
rect 12345 15311 12403 15317
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 5074 15104 5080 15156
rect 5132 15104 5138 15156
rect 6638 15104 6644 15156
rect 6696 15144 6702 15156
rect 9674 15144 9680 15156
rect 6696 15116 9680 15144
rect 6696 15104 6702 15116
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 11054 15144 11060 15156
rect 10735 15116 11060 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12345 15147 12403 15153
rect 12345 15144 12357 15147
rect 12308 15116 12357 15144
rect 12308 15104 12314 15116
rect 12345 15113 12357 15116
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 13446 15104 13452 15156
rect 13504 15144 13510 15156
rect 13541 15147 13599 15153
rect 13541 15144 13553 15147
rect 13504 15116 13553 15144
rect 13504 15104 13510 15116
rect 13541 15113 13553 15116
rect 13587 15113 13599 15147
rect 13541 15107 13599 15113
rect 6730 15036 6736 15088
rect 6788 15036 6794 15088
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 7190 15076 7196 15088
rect 6880 15048 7196 15076
rect 6880 15036 6886 15048
rect 7190 15036 7196 15048
rect 7248 15036 7254 15088
rect 7653 15011 7711 15017
rect 6472 14980 7328 15008
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14940 5319 14943
rect 5442 14940 5448 14952
rect 5307 14912 5448 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5442 14900 5448 14912
rect 5500 14900 5506 14952
rect 5626 14900 5632 14952
rect 5684 14940 5690 14952
rect 6472 14949 6500 14980
rect 6273 14943 6331 14949
rect 6273 14940 6285 14943
rect 5684 14912 6285 14940
rect 5684 14900 5690 14912
rect 6273 14909 6285 14912
rect 6319 14909 6331 14943
rect 6273 14903 6331 14909
rect 6457 14943 6515 14949
rect 6457 14909 6469 14943
rect 6503 14909 6515 14943
rect 6457 14903 6515 14909
rect 6549 14943 6607 14949
rect 6549 14909 6561 14943
rect 6595 14940 6607 14943
rect 6822 14940 6828 14952
rect 6595 14912 6828 14940
rect 6595 14909 6607 14912
rect 6549 14903 6607 14909
rect 6288 14872 6316 14903
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 6917 14875 6975 14881
rect 6917 14872 6929 14875
rect 6288 14844 6929 14872
rect 6564 14816 6592 14844
rect 6917 14841 6929 14844
rect 6963 14841 6975 14875
rect 7300 14872 7328 14980
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 7834 15008 7840 15020
rect 7699 14980 7840 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 14918 14968 14924 15020
rect 14976 14968 14982 15020
rect 7374 14900 7380 14952
rect 7432 14900 7438 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 8018 14940 8024 14952
rect 7515 14912 8024 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 10410 14900 10416 14952
rect 10468 14940 10474 14952
rect 10505 14943 10563 14949
rect 10505 14940 10517 14943
rect 10468 14912 10517 14940
rect 10468 14900 10474 14912
rect 10505 14909 10517 14912
rect 10551 14909 10563 14943
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 10505 14903 10563 14909
rect 12544 14912 12817 14940
rect 8570 14872 8576 14884
rect 6917 14835 6975 14841
rect 7024 14844 8576 14872
rect 6086 14764 6092 14816
rect 6144 14764 6150 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 7024 14813 7052 14844
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 12161 14875 12219 14881
rect 12161 14872 12173 14875
rect 10836 14844 12173 14872
rect 10836 14832 10842 14844
rect 12161 14841 12173 14844
rect 12207 14841 12219 14875
rect 12161 14835 12219 14841
rect 7009 14807 7067 14813
rect 7009 14773 7021 14807
rect 7055 14773 7067 14807
rect 7009 14767 7067 14773
rect 7101 14807 7159 14813
rect 7101 14773 7113 14807
rect 7147 14804 7159 14807
rect 7190 14804 7196 14816
rect 7147 14776 7196 14804
rect 7147 14773 7159 14776
rect 7101 14767 7159 14773
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7282 14764 7288 14816
rect 7340 14764 7346 14816
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 7653 14807 7711 14813
rect 7653 14804 7665 14807
rect 7432 14776 7665 14804
rect 7432 14764 7438 14776
rect 7653 14773 7665 14776
rect 7699 14773 7711 14807
rect 7653 14767 7711 14773
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 10796 14804 10824 14832
rect 8168 14776 10824 14804
rect 8168 14764 8174 14776
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 12544 14813 12572 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 14654 14875 14712 14881
rect 14654 14872 14666 14875
rect 13004 14844 14666 14872
rect 13004 14813 13032 14844
rect 14654 14841 14666 14844
rect 14700 14841 14712 14875
rect 14654 14835 14712 14841
rect 12361 14807 12419 14813
rect 12361 14804 12373 14807
rect 12124 14776 12373 14804
rect 12124 14764 12130 14776
rect 12361 14773 12373 14776
rect 12407 14773 12419 14807
rect 12361 14767 12419 14773
rect 12529 14807 12587 14813
rect 12529 14773 12541 14807
rect 12575 14773 12587 14807
rect 12529 14767 12587 14773
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14773 13047 14807
rect 12989 14767 13047 14773
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 6822 14600 6828 14612
rect 4212 14572 6828 14600
rect 4212 14560 4218 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 10321 14603 10379 14609
rect 8904 14572 9260 14600
rect 8904 14560 8910 14572
rect 5429 14535 5487 14541
rect 5429 14501 5441 14535
rect 5475 14532 5487 14535
rect 5629 14535 5687 14541
rect 5475 14504 5580 14532
rect 5475 14501 5487 14504
rect 5429 14495 5487 14501
rect 5442 14396 5448 14408
rect 5276 14368 5448 14396
rect 5276 14337 5304 14368
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 5552 14328 5580 14504
rect 5629 14501 5641 14535
rect 5675 14501 5687 14535
rect 5629 14495 5687 14501
rect 6196 14504 6500 14532
rect 5644 14396 5672 14495
rect 6196 14473 6224 14504
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14433 6331 14467
rect 6472 14464 6500 14504
rect 6546 14492 6552 14544
rect 6604 14532 6610 14544
rect 8864 14532 8892 14560
rect 9232 14541 9260 14572
rect 10321 14569 10333 14603
rect 10367 14569 10379 14603
rect 10321 14563 10379 14569
rect 6604 14504 8892 14532
rect 9017 14535 9075 14541
rect 6604 14492 6610 14504
rect 9017 14501 9029 14535
rect 9063 14532 9075 14535
rect 9217 14535 9275 14541
rect 9063 14504 9168 14532
rect 9063 14501 9075 14504
rect 9017 14495 9075 14501
rect 9140 14476 9168 14504
rect 9217 14501 9229 14535
rect 9263 14501 9275 14535
rect 9217 14495 9275 14501
rect 9769 14535 9827 14541
rect 9769 14501 9781 14535
rect 9815 14532 9827 14535
rect 10336 14532 10364 14563
rect 10410 14560 10416 14612
rect 10468 14560 10474 14612
rect 11333 14603 11391 14609
rect 11333 14569 11345 14603
rect 11379 14600 11391 14603
rect 12158 14600 12164 14612
rect 11379 14572 12164 14600
rect 11379 14569 11391 14572
rect 11333 14563 11391 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12250 14560 12256 14612
rect 12308 14560 12314 14612
rect 12544 14572 13216 14600
rect 10565 14535 10623 14541
rect 10565 14532 10577 14535
rect 9815 14504 10272 14532
rect 10336 14504 10577 14532
rect 9815 14501 9827 14504
rect 9769 14495 9827 14501
rect 6472 14436 8708 14464
rect 6273 14427 6331 14433
rect 5644 14368 6224 14396
rect 6196 14340 6224 14368
rect 5997 14331 6055 14337
rect 5997 14328 6009 14331
rect 5552 14300 6009 14328
rect 5261 14291 5319 14297
rect 5997 14297 6009 14300
rect 6043 14297 6055 14331
rect 5997 14291 6055 14297
rect 6178 14288 6184 14340
rect 6236 14288 6242 14340
rect 6288 14328 6316 14427
rect 6638 14356 6644 14408
rect 6696 14356 6702 14408
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6880 14368 7021 14396
rect 6880 14356 6886 14368
rect 7009 14365 7021 14368
rect 7055 14396 7067 14399
rect 8202 14396 8208 14408
rect 7055 14368 8208 14396
rect 7055 14365 7067 14368
rect 7009 14359 7067 14365
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 8680 14396 8708 14436
rect 8754 14424 8760 14476
rect 8812 14424 8818 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9950 14464 9956 14476
rect 9180 14436 9956 14464
rect 9180 14424 9186 14436
rect 9950 14424 9956 14436
rect 10008 14464 10014 14476
rect 10045 14467 10103 14473
rect 10045 14464 10057 14467
rect 10008 14436 10057 14464
rect 10008 14424 10014 14436
rect 10045 14433 10057 14436
rect 10091 14433 10103 14467
rect 10244 14464 10272 14504
rect 10565 14501 10577 14504
rect 10611 14501 10623 14535
rect 10565 14495 10623 14501
rect 10778 14492 10784 14544
rect 10836 14492 10842 14544
rect 11698 14492 11704 14544
rect 11756 14492 11762 14544
rect 11793 14535 11851 14541
rect 11793 14501 11805 14535
rect 11839 14532 11851 14535
rect 12544 14532 12572 14572
rect 11839 14504 12572 14532
rect 11839 14501 11851 14504
rect 11793 14495 11851 14501
rect 12544 14476 12572 14504
rect 12621 14535 12679 14541
rect 12621 14501 12633 14535
rect 12667 14532 12679 14535
rect 12973 14535 13031 14541
rect 12667 14504 12940 14532
rect 12667 14501 12679 14504
rect 12621 14495 12679 14501
rect 11146 14464 11152 14476
rect 10244 14436 11152 14464
rect 10045 14427 10103 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14433 11483 14467
rect 11425 14427 11483 14433
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12342 14464 12348 14476
rect 11931 14436 12348 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 9677 14399 9735 14405
rect 8680 14368 9628 14396
rect 6362 14328 6368 14340
rect 6288 14300 6368 14328
rect 6362 14288 6368 14300
rect 6420 14328 6426 14340
rect 8849 14331 8907 14337
rect 8849 14328 8861 14331
rect 6420 14300 8861 14328
rect 6420 14288 6426 14300
rect 8849 14297 8861 14300
rect 8895 14297 8907 14331
rect 9600 14328 9628 14368
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9766 14396 9772 14408
rect 9723 14368 9772 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 11054 14396 11060 14408
rect 10183 14368 11060 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10152 14328 10180 14359
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 9600 14300 10180 14328
rect 11164 14328 11192 14424
rect 11440 14396 11468 14427
rect 12342 14424 12348 14436
rect 12400 14424 12406 14476
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12526 14464 12532 14476
rect 12483 14436 12532 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 12912 14464 12940 14504
rect 12973 14501 12985 14535
rect 13019 14532 13031 14535
rect 13078 14532 13084 14544
rect 13019 14504 13084 14532
rect 13019 14501 13031 14504
rect 12973 14495 13031 14501
rect 13078 14492 13084 14504
rect 13136 14492 13142 14544
rect 13188 14541 13216 14572
rect 13173 14535 13231 14541
rect 13173 14501 13185 14535
rect 13219 14532 13231 14535
rect 13446 14532 13452 14544
rect 13219 14504 13452 14532
rect 13219 14501 13231 14504
rect 13173 14495 13231 14501
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 12912 14436 13032 14464
rect 13004 14408 13032 14436
rect 11440 14368 12848 14396
rect 12820 14340 12848 14368
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 11164 14300 12081 14328
rect 8849 14291 8907 14297
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 12069 14291 12127 14297
rect 12158 14288 12164 14340
rect 12216 14328 12222 14340
rect 12434 14328 12440 14340
rect 12216 14300 12440 14328
rect 12216 14288 12222 14300
rect 12434 14288 12440 14300
rect 12492 14328 12498 14340
rect 12710 14328 12716 14340
rect 12492 14300 12716 14328
rect 12492 14288 12498 14300
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 12802 14288 12808 14340
rect 12860 14288 12866 14340
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 6086 14260 6092 14272
rect 5491 14232 6092 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 6086 14220 6092 14232
rect 6144 14220 6150 14272
rect 6196 14260 6224 14288
rect 8110 14260 8116 14272
rect 6196 14232 8116 14260
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8570 14220 8576 14272
rect 8628 14260 8634 14272
rect 9033 14263 9091 14269
rect 9033 14260 9045 14263
rect 8628 14232 9045 14260
rect 8628 14220 8634 14232
rect 9033 14229 9045 14232
rect 9079 14260 9091 14263
rect 9306 14260 9312 14272
rect 9079 14232 9312 14260
rect 9079 14229 9091 14232
rect 9033 14223 9091 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 10597 14263 10655 14269
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10965 14263 11023 14269
rect 10965 14260 10977 14263
rect 10643 14232 10977 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10965 14229 10977 14232
rect 11011 14229 11023 14263
rect 10965 14223 11023 14229
rect 11514 14220 11520 14272
rect 11572 14220 11578 14272
rect 11698 14220 11704 14272
rect 11756 14260 11762 14272
rect 12986 14260 12992 14272
rect 11756 14232 12992 14260
rect 11756 14220 11762 14232
rect 12986 14220 12992 14232
rect 13044 14220 13050 14272
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7006 14056 7012 14068
rect 6871 14028 7012 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7156 14028 8401 14056
rect 7156 14016 7162 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 8956 14028 9628 14056
rect 5721 13991 5779 13997
rect 5721 13957 5733 13991
rect 5767 13988 5779 13991
rect 6730 13988 6736 14000
rect 5767 13960 6736 13988
rect 5767 13957 5779 13960
rect 5721 13951 5779 13957
rect 6196 13864 6224 13960
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 6362 13880 6368 13932
rect 6420 13880 6426 13932
rect 6457 13923 6515 13929
rect 6457 13889 6469 13923
rect 6503 13920 6515 13923
rect 7098 13920 7104 13932
rect 6503 13892 7104 13920
rect 6503 13889 6515 13892
rect 6457 13883 6515 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8202 13880 8208 13932
rect 8260 13880 8266 13932
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 4212 13824 4353 13852
rect 4212 13812 4218 13824
rect 4341 13821 4353 13824
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 4608 13855 4666 13861
rect 4608 13821 4620 13855
rect 4654 13852 4666 13855
rect 5997 13855 6055 13861
rect 5997 13852 6009 13855
rect 4654 13824 6009 13852
rect 4654 13821 4666 13824
rect 4608 13815 4666 13821
rect 5997 13821 6009 13824
rect 6043 13821 6055 13855
rect 5997 13815 6055 13821
rect 6178 13812 6184 13864
rect 6236 13812 6242 13864
rect 6546 13812 6552 13864
rect 6604 13812 6610 13864
rect 6733 13855 6791 13861
rect 6733 13821 6745 13855
rect 6779 13852 6791 13855
rect 8389 13855 8447 13861
rect 8389 13852 8401 13855
rect 6779 13824 7236 13852
rect 6779 13821 6791 13824
rect 6733 13815 6791 13821
rect 5626 13744 5632 13796
rect 5684 13784 5690 13796
rect 6748 13784 6776 13815
rect 5684 13756 6776 13784
rect 5684 13744 5690 13756
rect 7208 13716 7236 13824
rect 7300 13824 8401 13852
rect 7300 13796 7328 13824
rect 8389 13821 8401 13824
rect 8435 13821 8447 13855
rect 8389 13815 8447 13821
rect 8570 13812 8576 13864
rect 8628 13812 8634 13864
rect 8956 13861 8984 14028
rect 9122 13948 9128 14000
rect 9180 13948 9186 14000
rect 9600 13988 9628 14028
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10226 14056 10232 14068
rect 9824 14028 10232 14056
rect 9824 14016 9830 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12345 14059 12403 14065
rect 12345 14056 12357 14059
rect 12124 14028 12357 14056
rect 12124 14016 12130 14028
rect 12345 14025 12357 14028
rect 12391 14025 12403 14059
rect 12345 14019 12403 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12618 14056 12624 14068
rect 12492 14028 12624 14056
rect 12492 14016 12498 14028
rect 12618 14016 12624 14028
rect 12676 14056 12682 14068
rect 13078 14056 13084 14068
rect 12676 14028 13084 14056
rect 12676 14016 12682 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 11698 13988 11704 14000
rect 9600 13960 11704 13988
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 12526 13988 12532 14000
rect 11808 13960 12532 13988
rect 9140 13920 9168 13948
rect 9585 13923 9643 13929
rect 9140 13892 9260 13920
rect 8941 13855 8999 13861
rect 8941 13852 8953 13855
rect 8680 13824 8953 13852
rect 7282 13744 7288 13796
rect 7340 13744 7346 13796
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 7938 13787 7996 13793
rect 7938 13784 7950 13787
rect 7708 13756 7950 13784
rect 7708 13744 7714 13756
rect 7938 13753 7950 13756
rect 7984 13753 7996 13787
rect 8680 13784 8708 13824
rect 8941 13821 8953 13824
rect 8987 13821 8999 13855
rect 8941 13815 8999 13821
rect 9122 13812 9128 13864
rect 9180 13812 9186 13864
rect 9232 13861 9260 13892
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 9674 13920 9680 13932
rect 9631 13892 9680 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 11514 13920 11520 13932
rect 9876 13892 11520 13920
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13821 9275 13855
rect 9217 13815 9275 13821
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9876 13861 9904 13892
rect 11514 13880 11520 13892
rect 11572 13880 11578 13932
rect 11808 13929 11836 13960
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 13541 13991 13599 13997
rect 13541 13988 13553 13991
rect 12768 13960 13553 13988
rect 12768 13948 12774 13960
rect 11793 13923 11851 13929
rect 11793 13889 11805 13923
rect 11839 13889 11851 13923
rect 12802 13920 12808 13932
rect 11793 13883 11851 13889
rect 12084 13892 12808 13920
rect 12084 13861 12112 13892
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9600 13824 9873 13852
rect 9600 13796 9628 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 7938 13747 7996 13753
rect 8496 13756 8708 13784
rect 8496 13716 8524 13756
rect 9582 13744 9588 13796
rect 9640 13744 9646 13796
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 9950 13784 9956 13796
rect 9723 13756 9956 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 7208 13688 8524 13716
rect 8846 13676 8852 13728
rect 8904 13716 8910 13728
rect 10060 13716 10088 13815
rect 12158 13812 12164 13864
rect 12216 13812 12222 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12268 13824 12449 13852
rect 11698 13744 11704 13796
rect 11756 13744 11762 13796
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12268 13784 12296 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12710 13812 12716 13864
rect 12768 13812 12774 13864
rect 12912 13852 12940 13960
rect 13541 13957 13553 13960
rect 13587 13957 13599 13991
rect 13541 13951 13599 13957
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 12986 13852 12992 13864
rect 12912 13824 12992 13852
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 14654 13855 14712 13861
rect 14654 13852 14666 13855
rect 13219 13824 14666 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 14654 13821 14666 13824
rect 14700 13821 14712 13855
rect 14654 13815 14712 13821
rect 11848 13756 12296 13784
rect 11848 13744 11854 13756
rect 12526 13716 12532 13728
rect 8904 13688 12532 13716
rect 8904 13676 8910 13688
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 5997 13515 6055 13521
rect 5997 13481 6009 13515
rect 6043 13512 6055 13515
rect 6546 13512 6552 13524
rect 6043 13484 6552 13512
rect 6043 13481 6055 13484
rect 5997 13475 6055 13481
rect 6546 13472 6552 13484
rect 6604 13472 6610 13524
rect 7650 13472 7656 13524
rect 7708 13472 7714 13524
rect 7834 13472 7840 13524
rect 7892 13472 7898 13524
rect 8754 13472 8760 13524
rect 8812 13521 8818 13524
rect 8812 13515 8841 13521
rect 8829 13512 8841 13515
rect 9582 13512 9588 13524
rect 8829 13484 9588 13512
rect 8829 13481 8841 13484
rect 8812 13475 8841 13481
rect 8812 13472 8818 13475
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 11146 13472 11152 13524
rect 11204 13512 11210 13524
rect 12158 13512 12164 13524
rect 11204 13484 12164 13512
rect 11204 13472 11210 13484
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 12618 13472 12624 13524
rect 12676 13512 12682 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12676 13484 12725 13512
rect 12676 13472 12682 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 12802 13472 12808 13524
rect 12860 13472 12866 13524
rect 12986 13472 12992 13524
rect 13044 13472 13050 13524
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 8573 13447 8631 13453
rect 7064 13416 7512 13444
rect 7064 13404 7070 13416
rect 6178 13336 6184 13388
rect 6236 13336 6242 13388
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13345 6975 13379
rect 6917 13339 6975 13345
rect 6362 13268 6368 13320
rect 6420 13268 6426 13320
rect 6932 13240 6960 13339
rect 7098 13336 7104 13388
rect 7156 13336 7162 13388
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 7374 13376 7380 13388
rect 7239 13348 7380 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7484 13385 7512 13416
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 8619 13416 9076 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13376 7527 13379
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 7515 13348 7757 13376
rect 7515 13345 7527 13348
rect 7469 13339 7527 13345
rect 7745 13345 7757 13348
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 7926 13336 7932 13388
rect 7984 13336 7990 13388
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7374 13240 7380 13252
rect 6932 13212 7380 13240
rect 7374 13200 7380 13212
rect 7432 13240 7438 13252
rect 8110 13240 8116 13252
rect 7432 13212 8116 13240
rect 7432 13200 7438 13212
rect 8110 13200 8116 13212
rect 8168 13200 8174 13252
rect 9048 13249 9076 13416
rect 9674 13404 9680 13456
rect 9732 13444 9738 13456
rect 10146 13447 10204 13453
rect 10146 13444 10158 13447
rect 9732 13416 10158 13444
rect 9732 13404 9738 13416
rect 10146 13413 10158 13416
rect 10192 13413 10204 13447
rect 10146 13407 10204 13413
rect 11514 13404 11520 13456
rect 11572 13444 11578 13456
rect 12066 13444 12072 13456
rect 11572 13416 12072 13444
rect 11572 13404 11578 13416
rect 12066 13404 12072 13416
rect 12124 13444 12130 13456
rect 12820 13444 12848 13472
rect 12124 13416 12664 13444
rect 12820 13416 13124 13444
rect 12124 13404 12130 13416
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 10962 13376 10968 13388
rect 10459 13348 10968 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13345 12587 13379
rect 12636 13376 12664 13416
rect 13096 13385 13124 13416
rect 12805 13379 12863 13385
rect 12805 13376 12817 13379
rect 12636 13348 12817 13376
rect 12529 13339 12587 13345
rect 12805 13345 12817 13348
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 13081 13379 13139 13385
rect 13081 13345 13093 13379
rect 13127 13345 13139 13379
rect 13081 13339 13139 13345
rect 11698 13268 11704 13320
rect 11756 13308 11762 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 11756 13280 12357 13308
rect 11756 13268 11762 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12544 13308 12572 13339
rect 12986 13308 12992 13320
rect 12544 13280 12992 13308
rect 12345 13271 12403 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 9033 13243 9091 13249
rect 9033 13209 9045 13243
rect 9079 13240 9091 13243
rect 9306 13240 9312 13252
rect 9079 13212 9312 13240
rect 9079 13209 9091 13212
rect 9033 13203 9091 13209
rect 9306 13200 9312 13212
rect 9364 13200 9370 13252
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 12805 13243 12863 13249
rect 12805 13240 12817 13243
rect 12768 13212 12817 13240
rect 12768 13200 12774 13212
rect 12805 13209 12817 13212
rect 12851 13209 12863 13243
rect 12805 13203 12863 13209
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 8846 13172 8852 13184
rect 8803 13144 8852 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 6641 12971 6699 12977
rect 6641 12937 6653 12971
rect 6687 12968 6699 12971
rect 6822 12968 6828 12980
rect 6687 12940 6828 12968
rect 6687 12937 6699 12940
rect 6641 12931 6699 12937
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 9122 12928 9128 12980
rect 9180 12928 9186 12980
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9582 12968 9588 12980
rect 9364 12940 9588 12968
rect 9364 12928 9370 12940
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11514 12968 11520 12980
rect 11112 12940 11520 12968
rect 11112 12928 11118 12940
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 13078 12928 13084 12980
rect 13136 12968 13142 12980
rect 14921 12971 14979 12977
rect 14921 12968 14933 12971
rect 13136 12940 14933 12968
rect 13136 12928 13142 12940
rect 14921 12937 14933 12940
rect 14967 12937 14979 12971
rect 14921 12931 14979 12937
rect 10045 12903 10103 12909
rect 10045 12900 10057 12903
rect 9508 12872 10057 12900
rect 5721 12835 5779 12841
rect 5721 12832 5733 12835
rect 5276 12804 5733 12832
rect 5276 12773 5304 12804
rect 5721 12801 5733 12804
rect 5767 12801 5779 12835
rect 5721 12795 5779 12801
rect 6178 12792 6184 12844
rect 6236 12832 6242 12844
rect 6236 12804 6868 12832
rect 6236 12792 6242 12804
rect 5261 12767 5319 12773
rect 5261 12733 5273 12767
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 5445 12767 5503 12773
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 5534 12764 5540 12776
rect 5491 12736 5540 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 4982 12588 4988 12640
rect 5040 12588 5046 12640
rect 5368 12628 5396 12727
rect 5534 12724 5540 12736
rect 5592 12724 5598 12776
rect 5626 12724 5632 12776
rect 5684 12724 5690 12776
rect 6365 12767 6423 12773
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 6380 12696 6408 12727
rect 6454 12696 6460 12708
rect 6380 12668 6460 12696
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 6546 12628 6552 12640
rect 5368 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 6638 12588 6644 12640
rect 6696 12637 6702 12640
rect 6840 12637 6868 12804
rect 8938 12792 8944 12844
rect 8996 12832 9002 12844
rect 8996 12804 9444 12832
rect 8996 12792 9002 12804
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8570 12764 8576 12776
rect 8444 12736 8576 12764
rect 8444 12724 8450 12736
rect 8570 12724 8576 12736
rect 8628 12764 8634 12776
rect 9416 12773 9444 12804
rect 9309 12767 9367 12773
rect 9309 12764 9321 12767
rect 8628 12736 9321 12764
rect 8628 12724 8634 12736
rect 9309 12733 9321 12736
rect 9355 12733 9367 12767
rect 9309 12727 9367 12733
rect 9401 12767 9459 12773
rect 9401 12733 9413 12767
rect 9447 12733 9459 12767
rect 9401 12727 9459 12733
rect 9324 12696 9352 12727
rect 9508 12696 9536 12872
rect 10045 12869 10057 12872
rect 10091 12869 10103 12903
rect 11808 12900 11836 12928
rect 11808 12872 12112 12900
rect 10045 12863 10103 12869
rect 9582 12792 9588 12844
rect 9640 12832 9646 12844
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 9640 12804 9689 12832
rect 9640 12792 9646 12804
rect 9677 12801 9689 12804
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 11698 12792 11704 12844
rect 11756 12832 11762 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 11756 12804 11805 12832
rect 11756 12792 11762 12804
rect 11793 12801 11805 12804
rect 11839 12832 11851 12835
rect 11882 12832 11888 12844
rect 11839 12804 11888 12832
rect 11839 12801 11851 12804
rect 11793 12795 11851 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 10318 12764 10324 12776
rect 9907 12736 10324 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 10318 12724 10324 12736
rect 10376 12724 10382 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11333 12767 11391 12773
rect 11333 12764 11345 12767
rect 11204 12736 11345 12764
rect 11204 12724 11210 12736
rect 11333 12733 11345 12736
rect 11379 12733 11391 12767
rect 11333 12727 11391 12733
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12733 12035 12767
rect 12084 12764 12112 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 12584 12872 12664 12900
rect 12584 12860 12590 12872
rect 12636 12841 12664 12872
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12621 12835 12679 12841
rect 12207 12804 12480 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12452 12773 12480 12804
rect 12621 12801 12633 12835
rect 12667 12832 12679 12835
rect 12986 12832 12992 12844
rect 12667 12804 12992 12832
rect 12667 12801 12679 12804
rect 12621 12795 12679 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12084 12736 12265 12764
rect 11977 12727 12035 12733
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 9324 12668 9536 12696
rect 9769 12699 9827 12705
rect 9769 12665 9781 12699
rect 9815 12665 9827 12699
rect 11992 12696 12020 12727
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 12805 12767 12863 12773
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 13078 12764 13084 12776
rect 12851 12736 13084 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 12820 12696 12848 12727
rect 13078 12724 13084 12736
rect 13136 12724 13142 12776
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12764 13599 12767
rect 13587 12736 13952 12764
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 13924 12708 13952 12736
rect 11992 12668 12848 12696
rect 12989 12699 13047 12705
rect 9769 12659 9827 12665
rect 12989 12665 13001 12699
rect 13035 12696 13047 12699
rect 13786 12699 13844 12705
rect 13786 12696 13798 12699
rect 13035 12668 13798 12696
rect 13035 12665 13047 12668
rect 12989 12659 13047 12665
rect 13786 12665 13798 12668
rect 13832 12665 13844 12699
rect 13786 12659 13844 12665
rect 6696 12631 6715 12637
rect 6703 12597 6715 12631
rect 6696 12591 6715 12597
rect 6825 12631 6883 12637
rect 6825 12597 6837 12631
rect 6871 12628 6883 12631
rect 8846 12628 8852 12640
rect 6871 12600 8852 12628
rect 6871 12597 6883 12600
rect 6825 12591 6883 12597
rect 6696 12588 6702 12591
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 9784 12628 9812 12659
rect 13906 12656 13912 12708
rect 13964 12656 13970 12708
rect 9640 12600 9812 12628
rect 9640 12588 9646 12600
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5905 12427 5963 12433
rect 5905 12424 5917 12427
rect 5592 12396 5917 12424
rect 5592 12384 5598 12396
rect 5905 12393 5917 12396
rect 5951 12393 5963 12427
rect 5905 12387 5963 12393
rect 7190 12384 7196 12436
rect 7248 12384 7254 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7834 12424 7840 12436
rect 7432 12396 7840 12424
rect 7432 12384 7438 12396
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 7926 12384 7932 12436
rect 7984 12424 7990 12436
rect 9582 12424 9588 12436
rect 7984 12396 9588 12424
rect 7984 12384 7990 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10134 12384 10140 12436
rect 10192 12384 10198 12436
rect 12894 12424 12900 12436
rect 11072 12396 12900 12424
rect 4424 12359 4482 12365
rect 4424 12325 4436 12359
rect 4470 12356 4482 12359
rect 4982 12356 4988 12368
rect 4470 12328 4988 12356
rect 4470 12325 4482 12328
rect 4424 12319 4482 12325
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 6730 12316 6736 12368
rect 6788 12356 6794 12368
rect 6917 12359 6975 12365
rect 6917 12356 6929 12359
rect 6788 12328 6929 12356
rect 6788 12316 6794 12328
rect 6917 12325 6929 12328
rect 6963 12325 6975 12359
rect 6917 12319 6975 12325
rect 7009 12359 7067 12365
rect 7009 12325 7021 12359
rect 7055 12356 7067 12359
rect 8754 12356 8760 12368
rect 7055 12328 8760 12356
rect 7055 12325 7067 12328
rect 7009 12319 7067 12325
rect 8754 12316 8760 12328
rect 8812 12316 8818 12368
rect 10962 12356 10968 12368
rect 9508 12328 10968 12356
rect 4154 12248 4160 12300
rect 4212 12248 4218 12300
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 6822 12288 6828 12300
rect 6696 12260 6828 12288
rect 6696 12248 6702 12260
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6362 12220 6368 12232
rect 6135 12192 6368 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7576 12220 7604 12251
rect 7742 12248 7748 12300
rect 7800 12248 7806 12300
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12288 7895 12291
rect 8110 12288 8116 12300
rect 7883 12260 8116 12288
rect 7883 12257 7895 12260
rect 7837 12251 7895 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 9508 12288 9536 12328
rect 10962 12316 10968 12328
rect 11020 12316 11026 12368
rect 11072 12300 11100 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 12989 12427 13047 12433
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13078 12424 13084 12436
rect 13035 12396 13084 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13078 12384 13084 12396
rect 13136 12384 13142 12436
rect 12710 12316 12716 12368
rect 12768 12316 12774 12368
rect 8260 12260 9536 12288
rect 8260 12248 8266 12260
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9640 12260 9812 12288
rect 9640 12248 9646 12260
rect 8018 12220 8024 12232
rect 6595 12192 7512 12220
rect 7576 12192 8024 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 5537 12155 5595 12161
rect 5537 12121 5549 12155
rect 5583 12152 5595 12155
rect 6472 12152 6500 12180
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5583 12124 6653 12152
rect 5583 12121 5595 12124
rect 5537 12115 5595 12121
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 7484 12152 7512 12192
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9784 12229 9812 12260
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10318 12288 10324 12300
rect 9916 12260 10324 12288
rect 9916 12248 9922 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 11054 12248 11060 12300
rect 11112 12248 11118 12300
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12124 12260 12817 12288
rect 12124 12248 12130 12260
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 13078 12248 13084 12300
rect 13136 12248 13142 12300
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 9950 12220 9956 12232
rect 9815 12192 9956 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 7926 12152 7932 12164
rect 7484 12124 7932 12152
rect 6641 12115 6699 12121
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7432 12056 7573 12084
rect 7432 12044 7438 12056
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7561 12047 7619 12053
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8202 12084 8208 12096
rect 7800 12056 8208 12084
rect 7800 12044 7806 12056
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 9030 12044 9036 12096
rect 9088 12084 9094 12096
rect 9493 12087 9551 12093
rect 9493 12084 9505 12087
rect 9088 12056 9505 12084
rect 9088 12044 9094 12056
rect 9493 12053 9505 12056
rect 9539 12053 9551 12087
rect 9692 12084 9720 12183
rect 9950 12180 9956 12192
rect 10008 12180 10014 12232
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10505 12155 10563 12161
rect 10505 12152 10517 12155
rect 10192 12124 10517 12152
rect 10192 12112 10198 12124
rect 10505 12121 10517 12124
rect 10551 12152 10563 12155
rect 11146 12152 11152 12164
rect 10551 12124 11152 12152
rect 10551 12121 10563 12124
rect 10505 12115 10563 12121
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 12526 12112 12532 12164
rect 12584 12152 12590 12164
rect 12805 12155 12863 12161
rect 12805 12152 12817 12155
rect 12584 12124 12817 12152
rect 12584 12112 12590 12124
rect 12805 12121 12817 12124
rect 12851 12121 12863 12155
rect 12805 12115 12863 12121
rect 10870 12084 10876 12096
rect 9692 12056 10876 12084
rect 9493 12047 9551 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 5960 11852 6500 11880
rect 5960 11840 5966 11852
rect 5445 11815 5503 11821
rect 5445 11781 5457 11815
rect 5491 11812 5503 11815
rect 6472 11812 6500 11852
rect 8018 11840 8024 11892
rect 8076 11840 8082 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8389 11883 8447 11889
rect 8389 11880 8401 11883
rect 8168 11852 8401 11880
rect 8168 11840 8174 11852
rect 8389 11849 8401 11852
rect 8435 11849 8447 11883
rect 8389 11843 8447 11849
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 13630 11880 13636 11892
rect 8904 11852 13636 11880
rect 8904 11840 8910 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 5491 11784 6408 11812
rect 6472 11784 11560 11812
rect 5491 11781 5503 11784
rect 5445 11775 5503 11781
rect 6380 11753 6408 11784
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11676 4123 11679
rect 4154 11676 4160 11688
rect 4111 11648 4160 11676
rect 4111 11645 4123 11648
rect 4065 11639 4123 11645
rect 4154 11636 4160 11648
rect 4212 11636 4218 11688
rect 4332 11611 4390 11617
rect 4332 11577 4344 11611
rect 4378 11608 4390 11611
rect 5718 11608 5724 11620
rect 4378 11580 5724 11608
rect 4378 11577 4390 11580
rect 4332 11571 4390 11577
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 6380 11608 6408 11707
rect 6546 11704 6552 11756
rect 6604 11744 6610 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 6604 11716 7297 11744
rect 6604 11704 6610 11716
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 6840 11685 6868 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7285 11707 7343 11713
rect 7392 11716 7665 11744
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6512 11648 6745 11676
rect 6512 11636 6518 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11645 6883 11679
rect 7392 11676 7420 11716
rect 7653 11713 7665 11716
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7892 11716 7941 11744
rect 7892 11704 7898 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8846 11704 8852 11756
rect 8904 11704 8910 11756
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 8987 11716 9812 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 6825 11639 6883 11645
rect 7116 11648 7420 11676
rect 6638 11608 6644 11620
rect 6380 11580 6644 11608
rect 6638 11568 6644 11580
rect 6696 11608 6702 11620
rect 7116 11617 7144 11648
rect 7466 11636 7472 11688
rect 7524 11636 7530 11688
rect 8202 11636 8208 11688
rect 8260 11636 8266 11688
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9784 11676 9812 11716
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 9950 11704 9956 11756
rect 10008 11744 10014 11756
rect 11532 11753 11560 11784
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12124 11784 12296 11812
rect 12124 11772 12130 11784
rect 12268 11753 12296 11784
rect 11517 11747 11575 11753
rect 10008 11716 11468 11744
rect 10008 11704 10014 11716
rect 10226 11676 10232 11688
rect 9784 11648 10232 11676
rect 9585 11639 9643 11645
rect 7101 11611 7159 11617
rect 7101 11608 7113 11611
rect 6696 11580 7113 11608
rect 6696 11568 6702 11580
rect 7101 11577 7113 11580
rect 7147 11577 7159 11611
rect 7101 11571 7159 11577
rect 7193 11611 7251 11617
rect 7193 11577 7205 11611
rect 7239 11608 7251 11611
rect 7926 11608 7932 11620
rect 7239 11580 7932 11608
rect 7239 11577 7251 11580
rect 7193 11571 7251 11577
rect 7926 11568 7932 11580
rect 7984 11568 7990 11620
rect 9600 11608 9628 11639
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 11440 11685 11468 11716
rect 11517 11713 11529 11747
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11744 11759 11747
rect 12253 11747 12311 11753
rect 11747 11716 12112 11744
rect 11747 11713 11759 11716
rect 11701 11707 11759 11713
rect 11425 11679 11483 11685
rect 11425 11645 11437 11679
rect 11471 11676 11483 11679
rect 11606 11676 11612 11688
rect 11471 11648 11612 11676
rect 11471 11645 11483 11648
rect 11425 11639 11483 11645
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12084 11685 12112 11716
rect 12253 11713 12265 11747
rect 12299 11713 12311 11747
rect 15102 11744 15108 11756
rect 12253 11707 12311 11713
rect 12544 11716 15108 11744
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11716 11648 11897 11676
rect 11716 11620 11744 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12544 11676 12572 11716
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 12483 11648 12572 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 9858 11608 9864 11620
rect 9600 11580 9864 11608
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 9953 11611 10011 11617
rect 9953 11577 9965 11611
rect 9999 11608 10011 11611
rect 10778 11608 10784 11620
rect 9999 11580 10784 11608
rect 9999 11577 10011 11580
rect 9953 11571 10011 11577
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 11698 11568 11704 11620
rect 11756 11568 11762 11620
rect 5813 11543 5871 11549
rect 5813 11509 5825 11543
rect 5859 11540 5871 11543
rect 6086 11540 6092 11552
rect 5859 11512 6092 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6270 11500 6276 11552
rect 6328 11540 6334 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6328 11512 6561 11540
rect 6328 11500 6334 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6549 11503 6607 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7466 11540 7472 11552
rect 6788 11512 7472 11540
rect 6788 11500 6794 11512
rect 7466 11500 7472 11512
rect 7524 11500 7530 11552
rect 8754 11500 8760 11552
rect 8812 11500 8818 11552
rect 9585 11543 9643 11549
rect 9585 11509 9597 11543
rect 9631 11540 9643 11543
rect 9674 11540 9680 11552
rect 9631 11512 9680 11540
rect 9631 11509 9643 11512
rect 9585 11503 9643 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 10045 11543 10103 11549
rect 10045 11509 10057 11543
rect 10091 11540 10103 11543
rect 10318 11540 10324 11552
rect 10091 11512 10324 11540
rect 10091 11509 10103 11512
rect 10045 11503 10103 11509
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10962 11540 10968 11552
rect 10459 11512 10968 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 11146 11540 11152 11552
rect 11103 11512 11152 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 12544 11540 12572 11648
rect 12986 11636 12992 11688
rect 13044 11676 13050 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13044 11648 13737 11676
rect 13044 11636 13050 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 12621 11611 12679 11617
rect 12621 11577 12633 11611
rect 12667 11608 12679 11611
rect 13998 11608 14004 11620
rect 12667 11580 14004 11608
rect 12667 11577 12679 11580
rect 12621 11571 12679 11577
rect 13998 11568 14004 11580
rect 14056 11568 14062 11620
rect 11572 11512 12572 11540
rect 11572 11500 11578 11512
rect 13906 11500 13912 11552
rect 13964 11500 13970 11552
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 5813 11339 5871 11345
rect 5813 11336 5825 11339
rect 5776 11308 5825 11336
rect 5776 11296 5782 11308
rect 5813 11305 5825 11308
rect 5859 11305 5871 11339
rect 5813 11299 5871 11305
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 8386 11336 8392 11348
rect 6512 11308 8392 11336
rect 6512 11296 6518 11308
rect 8386 11296 8392 11308
rect 8444 11336 8450 11348
rect 9306 11336 9312 11348
rect 8444 11308 9312 11336
rect 8444 11296 8450 11308
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 10778 11296 10784 11348
rect 10836 11296 10842 11348
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12158 11336 12164 11348
rect 12115 11308 12164 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12986 11296 12992 11348
rect 13044 11296 13050 11348
rect 6362 11268 6368 11280
rect 6196 11240 6368 11268
rect 6086 11160 6092 11212
rect 6144 11160 6150 11212
rect 6196 11209 6224 11240
rect 6362 11228 6368 11240
rect 6420 11268 6426 11280
rect 6730 11268 6736 11280
rect 6420 11240 6736 11268
rect 6420 11228 6426 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7374 11228 7380 11280
rect 7432 11228 7438 11280
rect 10229 11271 10287 11277
rect 10229 11237 10241 11271
rect 10275 11268 10287 11271
rect 10594 11268 10600 11280
rect 10275 11240 10600 11268
rect 10275 11237 10287 11240
rect 10229 11231 10287 11237
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 10962 11228 10968 11280
rect 11020 11268 11026 11280
rect 11020 11240 12434 11268
rect 11020 11228 11026 11240
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 6270 11160 6276 11212
rect 6328 11160 6334 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11200 6515 11203
rect 6638 11200 6644 11212
rect 6503 11172 6644 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6638 11160 6644 11172
rect 6696 11160 6702 11212
rect 7392 11200 7420 11228
rect 7653 11203 7711 11209
rect 7653 11200 7665 11203
rect 7392 11172 7665 11200
rect 7653 11169 7665 11172
rect 7699 11169 7711 11203
rect 7653 11163 7711 11169
rect 10505 11203 10563 11209
rect 10505 11169 10517 11203
rect 10551 11200 10563 11203
rect 11054 11200 11060 11212
rect 10551 11172 11060 11200
rect 10551 11169 10563 11172
rect 10505 11163 10563 11169
rect 11054 11160 11060 11172
rect 11112 11160 11118 11212
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 11974 11200 11980 11212
rect 11664 11172 11980 11200
rect 11664 11160 11670 11172
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12161 11203 12219 11209
rect 12161 11169 12173 11203
rect 12207 11169 12219 11203
rect 12406 11200 12434 11240
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 13265 11271 13323 11277
rect 13265 11268 13277 11271
rect 12952 11240 13277 11268
rect 12952 11228 12958 11240
rect 13265 11237 13277 11240
rect 13311 11237 13323 11271
rect 13265 11231 13323 11237
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12406 11172 12817 11200
rect 12161 11163 12219 11169
rect 12805 11169 12817 11172
rect 12851 11169 12863 11203
rect 12805 11163 12863 11169
rect 4154 11092 4160 11144
rect 4212 11132 4218 11144
rect 7374 11132 7380 11144
rect 4212 11104 7380 11132
rect 4212 11092 4218 11104
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8754 11132 8760 11144
rect 8352 11104 8760 11132
rect 8352 11092 8358 11104
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 10226 11132 10232 11144
rect 10183 11104 10232 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10870 11132 10876 11144
rect 10643 11104 10876 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10870 11092 10876 11104
rect 10928 11132 10934 11144
rect 11425 11135 11483 11141
rect 11425 11132 11437 11135
rect 10928 11104 11437 11132
rect 10928 11092 10934 11104
rect 11425 11101 11437 11104
rect 11471 11101 11483 11135
rect 12176 11132 12204 11163
rect 11425 11095 11483 11101
rect 11900 11104 12204 11132
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 6638 11064 6644 11076
rect 5684 11036 6644 11064
rect 5684 11024 5690 11036
rect 6638 11024 6644 11036
rect 6696 11024 6702 11076
rect 11900 11073 11928 11104
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 11885 11067 11943 11073
rect 11885 11033 11897 11067
rect 11931 11033 11943 11067
rect 11885 11027 11943 11033
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14553 10999 14611 11005
rect 14553 10996 14565 10999
rect 13872 10968 14565 10996
rect 13872 10956 13878 10968
rect 14553 10965 14565 10968
rect 14599 10965 14611 10999
rect 14553 10959 14611 10965
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 10870 10752 10876 10804
rect 10928 10752 10934 10804
rect 11054 10752 11060 10804
rect 11112 10752 11118 10804
rect 7098 10684 7104 10736
rect 7156 10724 7162 10736
rect 7285 10727 7343 10733
rect 7285 10724 7297 10727
rect 7156 10696 7297 10724
rect 7156 10684 7162 10696
rect 7285 10693 7297 10696
rect 7331 10693 7343 10727
rect 7285 10687 7343 10693
rect 10520 10696 11284 10724
rect 8202 10656 8208 10668
rect 7300 10628 8208 10656
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7300 10597 7328 10628
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10520 10665 10548 10696
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10376 10628 10517 10656
rect 10376 10616 10382 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11054 10656 11060 10668
rect 11011 10628 11060 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11256 10656 11284 10696
rect 13817 10659 13875 10665
rect 11256 10628 13768 10656
rect 7009 10591 7067 10597
rect 7009 10588 7021 10591
rect 6880 10560 7021 10588
rect 6880 10548 6886 10560
rect 7009 10557 7021 10560
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7285 10591 7343 10597
rect 7285 10557 7297 10591
rect 7331 10557 7343 10591
rect 7285 10551 7343 10557
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 10226 10588 10232 10600
rect 7984 10560 10232 10588
rect 7984 10548 7990 10560
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 11256 10597 11284 10628
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10744 10560 11161 10588
rect 10744 10548 10750 10560
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11241 10591 11299 10597
rect 11241 10557 11253 10591
rect 11287 10557 11299 10591
rect 11241 10551 11299 10557
rect 11517 10591 11575 10597
rect 11517 10557 11529 10591
rect 11563 10588 11575 10591
rect 12618 10588 12624 10600
rect 11563 10560 12624 10588
rect 11563 10557 11575 10560
rect 11517 10551 11575 10557
rect 6564 10492 7788 10520
rect 6564 10464 6592 10492
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6546 10452 6552 10464
rect 6236 10424 6552 10452
rect 6236 10412 6242 10424
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 6730 10412 6736 10464
rect 6788 10452 6794 10464
rect 7101 10455 7159 10461
rect 7101 10452 7113 10455
rect 6788 10424 7113 10452
rect 6788 10412 6794 10424
rect 7101 10421 7113 10424
rect 7147 10421 7159 10455
rect 7760 10452 7788 10492
rect 7834 10480 7840 10532
rect 7892 10520 7898 10532
rect 11532 10520 11560 10551
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10557 13599 10591
rect 13740 10588 13768 10628
rect 13817 10625 13829 10659
rect 13863 10656 13875 10659
rect 13998 10656 14004 10668
rect 13863 10628 14004 10656
rect 13863 10625 13875 10628
rect 13817 10619 13875 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 15654 10588 15660 10600
rect 13740 10560 15660 10588
rect 13541 10551 13599 10557
rect 11882 10520 11888 10532
rect 7892 10492 11560 10520
rect 11624 10492 11888 10520
rect 7892 10480 7898 10492
rect 8021 10455 8079 10461
rect 8021 10452 8033 10455
rect 7760 10424 8033 10452
rect 7101 10415 7159 10421
rect 8021 10421 8033 10424
rect 8067 10452 8079 10455
rect 11624 10452 11652 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 8067 10424 11652 10452
rect 8067 10421 8079 10424
rect 8021 10415 8079 10421
rect 11698 10412 11704 10464
rect 11756 10412 11762 10464
rect 13556 10452 13584 10551
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 13814 10452 13820 10464
rect 13556 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 18598 10452 18604 10464
rect 15160 10424 18604 10452
rect 15160 10412 15166 10424
rect 18598 10412 18604 10424
rect 18656 10412 18662 10464
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 6299 10251 6357 10257
rect 5644 10220 6224 10248
rect 5429 10183 5487 10189
rect 5429 10149 5441 10183
rect 5475 10180 5487 10183
rect 5534 10180 5540 10192
rect 5475 10152 5540 10180
rect 5475 10149 5487 10152
rect 5429 10143 5487 10149
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5644 10189 5672 10220
rect 5629 10183 5687 10189
rect 5629 10149 5641 10183
rect 5675 10149 5687 10183
rect 5629 10143 5687 10149
rect 6086 10140 6092 10192
rect 6144 10140 6150 10192
rect 6196 10180 6224 10220
rect 6299 10217 6311 10251
rect 6345 10248 6357 10251
rect 6822 10248 6828 10260
rect 6345 10220 6828 10248
rect 6345 10217 6357 10220
rect 6299 10211 6357 10217
rect 6822 10208 6828 10220
rect 6880 10248 6886 10260
rect 6880 10220 9352 10248
rect 6880 10208 6886 10220
rect 6196 10152 7052 10180
rect 6730 10112 6736 10124
rect 6288 10084 6736 10112
rect 4982 9868 4988 9920
rect 5040 9908 5046 9920
rect 5261 9911 5319 9917
rect 5261 9908 5273 9911
rect 5040 9880 5273 9908
rect 5040 9868 5046 9880
rect 5261 9877 5273 9880
rect 5307 9877 5319 9911
rect 5261 9871 5319 9877
rect 5445 9911 5503 9917
rect 5445 9877 5457 9911
rect 5491 9908 5503 9911
rect 5810 9908 5816 9920
rect 5491 9880 5816 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5810 9868 5816 9880
rect 5868 9868 5874 9920
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6288 9917 6316 10084
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 7024 10044 7052 10152
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 7469 10183 7527 10189
rect 7469 10180 7481 10183
rect 7432 10152 7481 10180
rect 7432 10140 7438 10152
rect 7469 10149 7481 10152
rect 7515 10149 7527 10183
rect 7469 10143 7527 10149
rect 9214 10140 9220 10192
rect 9272 10140 9278 10192
rect 9324 10180 9352 10220
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9769 10251 9827 10257
rect 9769 10248 9781 10251
rect 9548 10220 9781 10248
rect 9548 10208 9554 10220
rect 9769 10217 9781 10220
rect 9815 10217 9827 10251
rect 9769 10211 9827 10217
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 12710 10208 12716 10260
rect 12768 10208 12774 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13281 10251 13339 10257
rect 13281 10248 13293 10251
rect 12860 10220 13293 10248
rect 12860 10208 12866 10220
rect 13281 10217 13293 10220
rect 13327 10217 13339 10251
rect 13281 10211 13339 10217
rect 13449 10251 13507 10257
rect 13449 10217 13461 10251
rect 13495 10217 13507 10251
rect 13449 10211 13507 10217
rect 12437 10183 12495 10189
rect 12437 10180 12449 10183
rect 9324 10152 12449 10180
rect 12437 10149 12449 10152
rect 12483 10180 12495 10183
rect 12526 10180 12532 10192
rect 12483 10152 12532 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12636 10180 12664 10208
rect 13081 10183 13139 10189
rect 13081 10180 13093 10183
rect 12636 10152 13093 10180
rect 13081 10149 13093 10152
rect 13127 10149 13139 10183
rect 13081 10143 13139 10149
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7926 10112 7932 10124
rect 7147 10084 7932 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10226 10112 10232 10124
rect 9723 10084 10232 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 10468 10084 10517 10112
rect 10468 10072 10474 10084
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 10505 10075 10563 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 12621 10115 12679 10121
rect 12621 10081 12633 10115
rect 12667 10112 12679 10115
rect 12710 10112 12716 10124
rect 12667 10084 12716 10112
rect 12667 10081 12679 10084
rect 12621 10075 12679 10081
rect 7834 10044 7840 10056
rect 7024 10016 7840 10044
rect 7834 10004 7840 10016
rect 7892 10004 7898 10056
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10044 10011 10047
rect 10336 10044 10364 10072
rect 10980 10044 11008 10075
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10081 12863 10115
rect 13464 10112 13492 10211
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 13464 10084 13553 10112
rect 12805 10075 12863 10081
rect 13541 10081 13553 10084
rect 13587 10081 13599 10115
rect 13541 10075 13599 10081
rect 9999 10016 11008 10044
rect 12820 10044 12848 10075
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 14369 10115 14427 10121
rect 14369 10112 14381 10115
rect 13964 10084 14381 10112
rect 13964 10072 13970 10084
rect 14369 10081 14381 10084
rect 14415 10081 14427 10115
rect 14369 10075 14427 10081
rect 13078 10044 13084 10056
rect 12820 10016 13084 10044
rect 9999 10013 10011 10016
rect 9953 10007 10011 10013
rect 10520 9988 10548 10016
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13872 10016 14105 10044
rect 13872 10004 13878 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 7282 9936 7288 9988
rect 7340 9976 7346 9988
rect 8018 9976 8024 9988
rect 7340 9948 8024 9976
rect 7340 9936 7346 9948
rect 8018 9936 8024 9948
rect 8076 9936 8082 9988
rect 10502 9936 10508 9988
rect 10560 9936 10566 9988
rect 12986 9936 12992 9988
rect 13044 9936 13050 9988
rect 6273 9911 6331 9917
rect 6273 9908 6285 9911
rect 6236 9880 6285 9908
rect 6236 9868 6242 9880
rect 6273 9877 6285 9880
rect 6319 9877 6331 9911
rect 6273 9871 6331 9877
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6457 9911 6515 9917
rect 6457 9908 6469 9911
rect 6420 9880 6469 9908
rect 6420 9868 6426 9880
rect 6457 9877 6469 9880
rect 6503 9877 6515 9911
rect 6457 9871 6515 9877
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 8996 9880 9321 9908
rect 8996 9868 9002 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9766 9868 9772 9920
rect 9824 9908 9830 9920
rect 10137 9911 10195 9917
rect 10137 9908 10149 9911
rect 9824 9880 10149 9908
rect 9824 9868 9830 9880
rect 10137 9877 10149 9880
rect 10183 9877 10195 9911
rect 10137 9871 10195 9877
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11238 9908 11244 9920
rect 11112 9880 11244 9908
rect 11112 9868 11118 9880
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 13262 9868 13268 9920
rect 13320 9868 13326 9920
rect 13725 9911 13783 9917
rect 13725 9877 13737 9911
rect 13771 9908 13783 9911
rect 14090 9908 14096 9920
rect 13771 9880 14096 9908
rect 13771 9877 13783 9880
rect 13725 9871 13783 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16114 9908 16120 9920
rect 15712 9880 16120 9908
rect 15712 9868 15718 9880
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 5813 9707 5871 9713
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6086 9704 6092 9716
rect 5859 9676 6092 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6086 9664 6092 9676
rect 6144 9664 6150 9716
rect 8665 9707 8723 9713
rect 8665 9673 8677 9707
rect 8711 9704 8723 9707
rect 9214 9704 9220 9716
rect 8711 9676 9220 9704
rect 8711 9673 8723 9676
rect 8665 9667 8723 9673
rect 9214 9664 9220 9676
rect 9272 9664 9278 9716
rect 10410 9664 10416 9716
rect 10468 9664 10474 9716
rect 10597 9707 10655 9713
rect 10597 9673 10609 9707
rect 10643 9704 10655 9707
rect 10686 9704 10692 9716
rect 10643 9676 10692 9704
rect 10643 9673 10655 9676
rect 10597 9667 10655 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 11885 9707 11943 9713
rect 11885 9673 11897 9707
rect 11931 9704 11943 9707
rect 11931 9676 12940 9704
rect 11931 9673 11943 9676
rect 11885 9667 11943 9673
rect 6178 9596 6184 9648
rect 6236 9636 6242 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6236 9608 6653 9636
rect 6236 9596 6242 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 9766 9636 9772 9648
rect 6641 9599 6699 9605
rect 9048 9608 9772 9636
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 4212 9540 4445 9568
rect 4212 9528 4218 9540
rect 4433 9537 4445 9540
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 9048 9577 9076 9608
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 9953 9639 10011 9645
rect 9953 9605 9965 9639
rect 9999 9636 10011 9639
rect 10965 9639 11023 9645
rect 10965 9636 10977 9639
rect 9999 9608 10977 9636
rect 9999 9605 10011 9608
rect 9953 9599 10011 9605
rect 10965 9605 10977 9608
rect 11011 9605 11023 9639
rect 10965 9599 11023 9605
rect 12802 9596 12808 9648
rect 12860 9596 12866 9648
rect 12912 9645 12940 9676
rect 12897 9639 12955 9645
rect 12897 9605 12909 9639
rect 12943 9605 12955 9639
rect 12897 9599 12955 9605
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9033 9531 9091 9537
rect 5997 9503 6055 9509
rect 5997 9469 6009 9503
rect 6043 9500 6055 9503
rect 6178 9500 6184 9512
rect 6043 9472 6184 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7432 9472 8033 9500
rect 7432 9460 7438 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 9048 9500 9076 9531
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 9180 9540 9413 9568
rect 9180 9528 9186 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 8021 9463 8079 9469
rect 8772 9472 9076 9500
rect 4700 9435 4758 9441
rect 4700 9401 4712 9435
rect 4746 9432 4758 9435
rect 4890 9432 4896 9444
rect 4746 9404 4896 9432
rect 4746 9401 4758 9404
rect 4700 9395 4758 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 6549 9435 6607 9441
rect 6549 9401 6561 9435
rect 6595 9432 6607 9435
rect 7190 9432 7196 9444
rect 6595 9404 7196 9432
rect 6595 9401 6607 9404
rect 6549 9395 6607 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 7754 9435 7812 9441
rect 7754 9432 7766 9435
rect 7524 9404 7766 9432
rect 7524 9392 7530 9404
rect 7754 9401 7766 9404
rect 7800 9401 7812 9435
rect 8481 9435 8539 9441
rect 8481 9432 8493 9435
rect 7754 9395 7812 9401
rect 8404 9404 8493 9432
rect 8404 9376 8432 9404
rect 8481 9401 8493 9404
rect 8527 9401 8539 9435
rect 8481 9395 8539 9401
rect 8686 9435 8744 9441
rect 8686 9401 8698 9435
rect 8732 9432 8744 9435
rect 8772 9432 8800 9472
rect 9306 9460 9312 9512
rect 9364 9460 9370 9512
rect 9416 9500 9444 9531
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 9640 9540 10149 9568
rect 9640 9528 9646 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10594 9568 10600 9580
rect 10284 9540 10600 9568
rect 10284 9528 10290 9540
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 11882 9528 11888 9580
rect 11940 9568 11946 9580
rect 12158 9568 12164 9580
rect 11940 9540 12164 9568
rect 11940 9528 11946 9540
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12400 9540 12633 9568
rect 12400 9528 12406 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12768 9540 13400 9568
rect 12768 9528 12774 9540
rect 10045 9503 10103 9509
rect 10045 9500 10057 9503
rect 9416 9472 10057 9500
rect 10045 9469 10057 9472
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 8732 9404 8800 9432
rect 9677 9435 9735 9441
rect 8732 9401 8744 9404
rect 8686 9395 8744 9401
rect 9677 9401 9689 9435
rect 9723 9432 9735 9435
rect 9858 9432 9864 9444
rect 9723 9404 9864 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 10244 9441 10272 9528
rect 13372 9512 13400 9540
rect 10410 9460 10416 9512
rect 10468 9460 10474 9512
rect 10686 9460 10692 9512
rect 10744 9460 10750 9512
rect 12434 9500 12440 9512
rect 11716 9472 12440 9500
rect 10229 9435 10287 9441
rect 10229 9401 10241 9435
rect 10275 9401 10287 9435
rect 10428 9432 10456 9460
rect 10870 9432 10876 9444
rect 10428 9404 10876 9432
rect 10229 9395 10287 9401
rect 10870 9392 10876 9404
rect 10928 9432 10934 9444
rect 11716 9441 11744 9472
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12526 9460 12532 9512
rect 12584 9460 12590 9512
rect 13078 9460 13084 9512
rect 13136 9509 13142 9512
rect 13136 9503 13185 9509
rect 13136 9469 13139 9503
rect 13173 9500 13185 9503
rect 13173 9472 13308 9500
rect 13173 9469 13185 9472
rect 13136 9463 13185 9469
rect 13136 9460 13142 9463
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10928 9404 10977 9432
rect 10928 9392 10934 9404
rect 10965 9401 10977 9404
rect 11011 9401 11023 9435
rect 10965 9395 11023 9401
rect 11701 9435 11759 9441
rect 11701 9401 11713 9435
rect 11747 9401 11759 9435
rect 11701 9395 11759 9401
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12986 9432 12992 9444
rect 12299 9404 12992 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12986 9392 12992 9404
rect 13044 9392 13050 9444
rect 13280 9432 13308 9472
rect 13354 9460 13360 9512
rect 13412 9460 13418 9512
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 13280 9404 13400 9432
rect 6454 9324 6460 9376
rect 6512 9364 6518 9376
rect 8386 9364 8392 9376
rect 6512 9336 8392 9364
rect 6512 9324 6518 9336
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8846 9324 8852 9376
rect 8904 9324 8910 9376
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 9398 9324 9404 9376
rect 9456 9364 9462 9376
rect 9585 9367 9643 9373
rect 9585 9364 9597 9367
rect 9456 9336 9597 9364
rect 9456 9324 9462 9336
rect 9585 9333 9597 9336
rect 9631 9333 9643 9367
rect 9585 9327 9643 9333
rect 9766 9324 9772 9376
rect 9824 9324 9830 9376
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10429 9367 10487 9373
rect 10429 9364 10441 9367
rect 10376 9336 10441 9364
rect 10376 9324 10382 9336
rect 10429 9333 10441 9336
rect 10475 9333 10487 9367
rect 10429 9327 10487 9333
rect 10778 9324 10784 9376
rect 10836 9324 10842 9376
rect 11882 9324 11888 9376
rect 11940 9373 11946 9376
rect 11940 9367 11959 9373
rect 11947 9333 11959 9367
rect 11940 9327 11959 9333
rect 11940 9324 11946 9327
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 12952 9336 13277 9364
rect 12952 9324 12958 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13372 9364 13400 9404
rect 13814 9392 13820 9444
rect 13872 9432 13878 9444
rect 13970 9435 14028 9441
rect 13970 9432 13982 9435
rect 13872 9404 13982 9432
rect 13872 9392 13878 9404
rect 13970 9401 13982 9404
rect 14016 9401 14028 9435
rect 13970 9395 14028 9401
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 13372 9336 15117 9364
rect 13265 9327 13323 9333
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 4890 9120 4896 9172
rect 4948 9160 4954 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4948 9132 4997 9160
rect 4948 9120 4954 9132
rect 4985 9129 4997 9132
rect 5031 9129 5043 9163
rect 4985 9123 5043 9129
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 5905 9163 5963 9169
rect 5905 9160 5917 9163
rect 5592 9132 5917 9160
rect 5592 9120 5598 9132
rect 5905 9129 5917 9132
rect 5951 9129 5963 9163
rect 5905 9123 5963 9129
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7466 9160 7472 9172
rect 7423 9132 7472 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 9214 9120 9220 9172
rect 9272 9160 9278 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 9272 9132 9965 9160
rect 9272 9120 9278 9132
rect 9953 9129 9965 9132
rect 9999 9160 10011 9163
rect 10686 9160 10692 9172
rect 9999 9132 10692 9160
rect 9999 9129 10011 9132
rect 9953 9123 10011 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11940 9132 12173 9160
rect 11940 9120 11946 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 12161 9123 12219 9129
rect 13262 9120 13268 9172
rect 13320 9160 13326 9172
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 13320 9132 13461 9160
rect 13320 9120 13326 9132
rect 13449 9129 13461 9132
rect 13495 9129 13507 9163
rect 13449 9123 13507 9129
rect 13725 9163 13783 9169
rect 13725 9129 13737 9163
rect 13771 9160 13783 9163
rect 13814 9160 13820 9172
rect 13771 9132 13820 9160
rect 13771 9129 13783 9132
rect 13725 9123 13783 9129
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 6457 9095 6515 9101
rect 6457 9092 6469 9095
rect 6144 9064 6469 9092
rect 6144 9052 6150 9064
rect 6457 9061 6469 9064
rect 6503 9061 6515 9095
rect 6457 9055 6515 9061
rect 6546 9052 6552 9104
rect 6604 9052 6610 9104
rect 6914 9092 6920 9104
rect 6840 9064 6920 9092
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5169 9027 5227 9033
rect 5169 9024 5181 9027
rect 5040 8996 5181 9024
rect 5040 8984 5046 8996
rect 5169 8993 5181 8996
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 6181 9027 6239 9033
rect 6181 8993 6193 9027
rect 6227 9024 6239 9027
rect 6362 9024 6368 9036
rect 6227 8996 6368 9024
rect 6227 8993 6239 8996
rect 6181 8987 6239 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 6641 9027 6699 9033
rect 6641 8993 6653 9027
rect 6687 9024 6699 9027
rect 6730 9024 6736 9036
rect 6687 8996 6736 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6840 9033 6868 9064
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 8846 9052 8852 9104
rect 8904 9092 8910 9104
rect 10137 9095 10195 9101
rect 8904 9064 9628 9092
rect 8904 9052 8910 9064
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 7098 9024 7104 9036
rect 6825 8987 6883 8993
rect 6932 8996 7104 9024
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6454 8956 6460 8968
rect 6135 8928 6460 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6932 8965 6960 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 7190 8984 7196 9036
rect 7248 8984 7254 9036
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 9122 9024 9128 9036
rect 8076 8996 9128 9024
rect 8076 8984 8082 8996
rect 9122 8984 9128 8996
rect 9180 9024 9186 9036
rect 9306 9024 9312 9036
rect 9180 8996 9312 9024
rect 9180 8984 9186 8996
rect 9306 8984 9312 8996
rect 9364 8984 9370 9036
rect 9398 8984 9404 9036
rect 9456 8984 9462 9036
rect 9600 9024 9628 9064
rect 10137 9061 10149 9095
rect 10183 9092 10195 9095
rect 10502 9092 10508 9104
rect 10183 9064 10508 9092
rect 10183 9061 10195 9064
rect 10137 9055 10195 9061
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 14090 9101 14096 9104
rect 14084 9092 14096 9101
rect 12124 9064 13584 9092
rect 14051 9064 14096 9092
rect 12124 9052 12130 9064
rect 9674 9024 9680 9036
rect 9600 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9858 8984 9864 9036
rect 9916 8984 9922 9036
rect 10226 8984 10232 9036
rect 10284 9024 10290 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 10284 8996 10333 9024
rect 10284 8984 10290 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 9024 12495 9027
rect 12618 9024 12624 9036
rect 12483 8996 12624 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12710 8984 12716 9036
rect 12768 9024 12774 9036
rect 13078 9024 13084 9036
rect 12768 8996 13084 9024
rect 12768 8984 12774 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13354 9024 13360 9036
rect 13311 8996 13360 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13354 8984 13360 8996
rect 13412 8984 13418 9036
rect 13556 9033 13584 9064
rect 14084 9055 14096 9064
rect 14090 9052 14096 9055
rect 14148 9052 14154 9104
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 8993 13599 9027
rect 13541 8987 13599 8993
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8925 6975 8959
rect 6917 8919 6975 8925
rect 7009 8959 7067 8965
rect 7009 8925 7021 8959
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 6822 8888 6828 8900
rect 6328 8860 6828 8888
rect 6328 8848 6334 8860
rect 6822 8848 6828 8860
rect 6880 8888 6886 8900
rect 7024 8888 7052 8919
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 11146 8956 11152 8968
rect 8444 8928 11152 8956
rect 8444 8916 8450 8928
rect 11146 8916 11152 8928
rect 11204 8956 11210 8968
rect 12342 8956 12348 8968
rect 11204 8928 12348 8956
rect 11204 8916 11210 8928
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 6880 8860 7052 8888
rect 6880 8848 6886 8860
rect 12158 8848 12164 8900
rect 12216 8888 12222 8900
rect 12820 8888 12848 8919
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 13173 8959 13231 8965
rect 13173 8925 13185 8959
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 12216 8860 12848 8888
rect 12216 8848 12222 8860
rect 9214 8780 9220 8832
rect 9272 8780 9278 8832
rect 13004 8820 13032 8916
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 13188 8888 13216 8919
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13817 8959 13875 8965
rect 13817 8956 13829 8959
rect 13780 8928 13829 8956
rect 13780 8916 13786 8928
rect 13817 8925 13829 8928
rect 13863 8925 13875 8959
rect 13817 8919 13875 8925
rect 13136 8860 13216 8888
rect 13136 8848 13142 8860
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 13004 8792 15209 8820
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 15197 8783 15255 8789
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 5810 8576 5816 8628
rect 5868 8576 5874 8628
rect 7650 8616 7656 8628
rect 6564 8588 7656 8616
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8412 6055 8415
rect 6086 8412 6092 8424
rect 6043 8384 6092 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 6178 8372 6184 8424
rect 6236 8372 6242 8424
rect 6270 8372 6276 8424
rect 6328 8372 6334 8424
rect 6564 8421 6592 8588
rect 7650 8576 7656 8588
rect 7708 8616 7714 8628
rect 9490 8616 9496 8628
rect 7708 8588 9496 8616
rect 7708 8576 7714 8588
rect 9490 8576 9496 8588
rect 9548 8616 9554 8628
rect 9674 8616 9680 8628
rect 9548 8588 9680 8616
rect 9548 8576 9554 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 9916 8588 10333 8616
rect 9916 8576 9922 8588
rect 10321 8585 10333 8588
rect 10367 8585 10379 8619
rect 10321 8579 10379 8585
rect 12526 8576 12532 8628
rect 12584 8616 12590 8628
rect 12894 8616 12900 8628
rect 12584 8588 12900 8616
rect 12584 8576 12590 8588
rect 12894 8576 12900 8588
rect 12952 8616 12958 8628
rect 13078 8616 13084 8628
rect 12952 8588 13084 8616
rect 12952 8576 12958 8588
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 9692 8548 9720 8576
rect 10778 8548 10784 8560
rect 9692 8520 10784 8548
rect 10778 8508 10784 8520
rect 10836 8508 10842 8560
rect 12345 8551 12403 8557
rect 12345 8517 12357 8551
rect 12391 8548 12403 8551
rect 12618 8548 12624 8560
rect 12391 8520 12624 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 12618 8508 12624 8520
rect 12676 8508 12682 8560
rect 9306 8440 9312 8492
rect 9364 8480 9370 8492
rect 9364 8452 11284 8480
rect 9364 8440 9370 8452
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6638 8372 6644 8424
rect 6696 8412 6702 8424
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 6696 8384 6745 8412
rect 6696 8372 6702 8384
rect 6733 8381 6745 8384
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 6825 8415 6883 8421
rect 6825 8381 6837 8415
rect 6871 8412 6883 8415
rect 7282 8412 7288 8424
rect 6871 8384 7288 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 6748 8344 6776 8375
rect 7282 8372 7288 8384
rect 7340 8372 7346 8424
rect 8754 8372 8760 8424
rect 8812 8372 8818 8424
rect 8938 8372 8944 8424
rect 8996 8372 9002 8424
rect 9122 8372 9128 8424
rect 9180 8412 9186 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 9180 8384 9229 8412
rect 9180 8372 9186 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 10873 8415 10931 8421
rect 10873 8412 10885 8415
rect 10744 8384 10885 8412
rect 10744 8372 10750 8384
rect 10873 8381 10885 8384
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 11054 8372 11060 8424
rect 11112 8372 11118 8424
rect 11256 8421 11284 8452
rect 11241 8415 11299 8421
rect 11241 8381 11253 8415
rect 11287 8381 11299 8415
rect 11241 8375 11299 8381
rect 8294 8344 8300 8356
rect 6748 8316 8300 8344
rect 8294 8304 8300 8316
rect 8352 8304 8358 8356
rect 9306 8344 9312 8356
rect 9048 8316 9312 8344
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6328 8248 6377 8276
rect 6328 8236 6334 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6365 8239 6423 8245
rect 6730 8236 6736 8288
rect 6788 8276 6794 8288
rect 9048 8276 9076 8316
rect 9306 8304 9312 8316
rect 9364 8304 9370 8356
rect 12710 8304 12716 8356
rect 12768 8304 12774 8356
rect 6788 8248 9076 8276
rect 6788 8236 6794 8248
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9401 8279 9459 8285
rect 9401 8276 9413 8279
rect 9180 8248 9413 8276
rect 9180 8236 9186 8248
rect 9401 8245 9413 8248
rect 9447 8245 9459 8279
rect 9401 8239 9459 8245
rect 11146 8236 11152 8288
rect 11204 8236 11210 8288
rect 12513 8279 12571 8285
rect 12513 8245 12525 8279
rect 12559 8276 12571 8279
rect 13354 8276 13360 8288
rect 12559 8248 13360 8276
rect 12559 8245 12571 8248
rect 12513 8239 12571 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 8404 8044 9965 8072
rect 8404 8013 8432 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 9953 8035 10011 8041
rect 10965 8075 11023 8081
rect 10965 8041 10977 8075
rect 11011 8072 11023 8075
rect 11054 8072 11060 8084
rect 11011 8044 11060 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11330 8032 11336 8084
rect 11388 8032 11394 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12124 8044 12940 8072
rect 12124 8032 12130 8044
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 7973 8447 8007
rect 9769 8007 9827 8013
rect 8389 7967 8447 7973
rect 8772 7976 9444 8004
rect 8772 7948 8800 7976
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6012 7800 6040 7899
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6503 7908 6561 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7936 7619 7939
rect 7607 7908 8156 7936
rect 7607 7905 7619 7908
rect 7561 7899 7619 7905
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6012 7772 7297 7800
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7484 7800 7512 7831
rect 7650 7828 7656 7880
rect 7708 7828 7714 7880
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7868 7803 7871
rect 8018 7868 8024 7880
rect 7791 7840 8024 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8128 7868 8156 7908
rect 8202 7896 8208 7948
rect 8260 7936 8266 7948
rect 8297 7939 8355 7945
rect 8297 7936 8309 7939
rect 8260 7908 8309 7936
rect 8260 7896 8266 7908
rect 8297 7905 8309 7908
rect 8343 7936 8355 7939
rect 8343 7908 8708 7936
rect 8343 7905 8355 7908
rect 8297 7899 8355 7905
rect 8570 7868 8576 7880
rect 8128 7840 8576 7868
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 8680 7868 8708 7908
rect 8754 7896 8760 7948
rect 8812 7896 8818 7948
rect 9030 7896 9036 7948
rect 9088 7896 9094 7948
rect 9122 7896 9128 7948
rect 9180 7896 9186 7948
rect 9306 7896 9312 7948
rect 9364 7896 9370 7948
rect 9416 7945 9444 7976
rect 9769 7973 9781 8007
rect 9815 8004 9827 8007
rect 10226 8004 10232 8016
rect 9815 7976 10232 8004
rect 9815 7973 9827 7976
rect 9769 7967 9827 7973
rect 10226 7964 10232 7976
rect 10284 7964 10290 8016
rect 10321 8007 10379 8013
rect 10321 7973 10333 8007
rect 10367 8004 10379 8007
rect 11348 8004 11376 8032
rect 12526 8004 12532 8016
rect 10367 7976 11376 8004
rect 12176 7976 12532 8004
rect 10367 7973 10379 7976
rect 10321 7967 10379 7973
rect 9401 7939 9459 7945
rect 9401 7905 9413 7939
rect 9447 7905 9459 7939
rect 9401 7899 9459 7905
rect 9490 7896 9496 7948
rect 9548 7936 9554 7948
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 9548 7908 9597 7936
rect 9548 7896 9554 7908
rect 9585 7905 9597 7908
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 8846 7868 8852 7880
rect 8680 7840 8852 7868
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 9600 7868 9628 7899
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 10836 7908 11345 7936
rect 10836 7896 10842 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11974 7896 11980 7948
rect 12032 7896 12038 7948
rect 12176 7945 12204 7976
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7905 12219 7939
rect 12161 7899 12219 7905
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12713 7939 12771 7945
rect 12483 7908 12517 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12713 7905 12725 7939
rect 12759 7936 12771 7939
rect 12802 7936 12808 7948
rect 12759 7908 12808 7936
rect 12759 7905 12771 7908
rect 12713 7899 12771 7905
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 9600 7840 10425 7868
rect 8941 7831 8999 7837
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 10413 7831 10471 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 11238 7868 11244 7880
rect 10643 7840 11244 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 11238 7828 11244 7840
rect 11296 7868 11302 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11296 7840 11437 7868
rect 11296 7828 11302 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 12452 7868 12480 7899
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 12912 7945 12940 8044
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13170 7936 13176 7948
rect 13127 7908 13176 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13170 7896 13176 7908
rect 13228 7896 13234 7948
rect 13354 7868 13360 7880
rect 11517 7831 11575 7837
rect 12084 7840 13360 7868
rect 7484 7772 10732 7800
rect 7285 7763 7343 7769
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 6270 7732 6276 7744
rect 5859 7704 6276 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7834 7692 7840 7744
rect 7892 7732 7898 7744
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7892 7704 7941 7732
rect 7892 7692 7898 7704
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 7929 7695 7987 7701
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 8478 7732 8484 7744
rect 8159 7704 8484 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 8573 7735 8631 7741
rect 8573 7701 8585 7735
rect 8619 7732 8631 7735
rect 8662 7732 8668 7744
rect 8619 7704 8668 7732
rect 8619 7701 8631 7704
rect 8573 7695 8631 7701
rect 8662 7692 8668 7704
rect 8720 7692 8726 7744
rect 8938 7692 8944 7744
rect 8996 7732 9002 7744
rect 9490 7732 9496 7744
rect 8996 7704 9496 7732
rect 8996 7692 9002 7704
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10704 7732 10732 7772
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 11532 7800 11560 7831
rect 12084 7800 12112 7840
rect 12989 7803 13047 7809
rect 12989 7800 13001 7803
rect 11020 7772 12112 7800
rect 12176 7772 13001 7800
rect 11020 7760 11026 7772
rect 12176 7732 12204 7772
rect 12989 7769 13001 7772
rect 13035 7769 13047 7803
rect 12989 7763 13047 7769
rect 10704 7704 12204 7732
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12618 7732 12624 7744
rect 12391 7704 12624 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12710 7692 12716 7744
rect 12768 7692 12774 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 13096 7732 13124 7840
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 12952 7704 13124 7732
rect 12952 7692 12958 7704
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 6822 7528 6828 7540
rect 6604 7500 6828 7528
rect 6604 7488 6610 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 8570 7528 8576 7540
rect 7147 7500 8576 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 10962 7488 10968 7540
rect 11020 7488 11026 7540
rect 6270 7352 6276 7404
rect 6328 7352 6334 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 7374 7392 7380 7404
rect 6595 7364 7380 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 7374 7352 7380 7364
rect 7432 7392 7438 7404
rect 8110 7392 8116 7404
rect 7432 7364 8116 7392
rect 7432 7352 7438 7364
rect 8110 7352 8116 7364
rect 8168 7392 8174 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8168 7364 8401 7392
rect 8168 7352 8174 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 8846 7352 8852 7404
rect 8904 7392 8910 7404
rect 12345 7395 12403 7401
rect 8904 7364 9904 7392
rect 8904 7352 8910 7364
rect 6638 7284 6644 7336
rect 6696 7284 6702 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6880 7296 6929 7324
rect 6880 7284 6886 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 3694 7216 3700 7268
rect 3752 7256 3758 7268
rect 4893 7259 4951 7265
rect 4893 7256 4905 7259
rect 3752 7228 4905 7256
rect 3752 7216 3758 7228
rect 4893 7225 4905 7228
rect 4939 7225 4951 7259
rect 4893 7219 4951 7225
rect 4908 7188 4936 7219
rect 6546 7216 6552 7268
rect 6604 7256 6610 7268
rect 7300 7256 7328 7287
rect 8386 7256 8392 7268
rect 6604 7228 7328 7256
rect 7852 7228 8392 7256
rect 6604 7216 6610 7228
rect 6733 7191 6791 7197
rect 6733 7188 6745 7191
rect 4908 7160 6745 7188
rect 6733 7157 6745 7160
rect 6779 7188 6791 7191
rect 7098 7188 7104 7200
rect 6779 7160 7104 7188
rect 6779 7157 6791 7160
rect 6733 7151 6791 7157
rect 7098 7148 7104 7160
rect 7156 7188 7162 7200
rect 7852 7188 7880 7228
rect 8386 7216 8392 7228
rect 8444 7216 8450 7268
rect 7156 7160 7880 7188
rect 7929 7191 7987 7197
rect 7156 7148 7162 7160
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 8662 7188 8668 7200
rect 7975 7160 8668 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8662 7148 8668 7160
rect 8720 7148 8726 7200
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9769 7191 9827 7197
rect 9769 7188 9781 7191
rect 8812 7160 9781 7188
rect 8812 7148 8818 7160
rect 9769 7157 9781 7160
rect 9815 7157 9827 7191
rect 9876 7188 9904 7364
rect 12345 7361 12357 7395
rect 12391 7392 12403 7395
rect 13722 7392 13728 7404
rect 12391 7364 13728 7392
rect 12391 7361 12403 7364
rect 12345 7355 12403 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 12078 7327 12136 7333
rect 12078 7324 12090 7327
rect 11204 7296 12090 7324
rect 11204 7284 11210 7296
rect 12078 7293 12090 7296
rect 12124 7293 12136 7327
rect 12078 7287 12136 7293
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 11698 7216 11704 7268
rect 11756 7256 11762 7268
rect 12452 7256 12480 7287
rect 12618 7284 12624 7336
rect 12676 7284 12682 7336
rect 12710 7284 12716 7336
rect 12768 7284 12774 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 12894 7324 12900 7336
rect 12851 7296 12900 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 12989 7287 13047 7293
rect 11756 7228 12480 7256
rect 11756 7216 11762 7228
rect 12526 7216 12532 7268
rect 12584 7256 12590 7268
rect 13004 7256 13032 7287
rect 12584 7228 13032 7256
rect 12584 7216 12590 7228
rect 12802 7188 12808 7200
rect 9876 7160 12808 7188
rect 9769 7151 9827 7157
rect 12802 7148 12808 7160
rect 12860 7148 12866 7200
rect 13170 7148 13176 7200
rect 13228 7148 13234 7200
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 8849 6987 8907 6993
rect 6604 6956 8248 6984
rect 6604 6944 6610 6956
rect 8220 6925 8248 6956
rect 8849 6953 8861 6987
rect 8895 6984 8907 6987
rect 9674 6984 9680 6996
rect 8895 6956 9680 6984
rect 8895 6953 8907 6956
rect 8849 6947 8907 6953
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 12526 6984 12532 6996
rect 12391 6956 12532 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 8205 6919 8263 6925
rect 8205 6885 8217 6919
rect 8251 6885 8263 6919
rect 8405 6919 8463 6925
rect 8405 6916 8417 6919
rect 8205 6879 8263 6885
rect 8404 6885 8417 6916
rect 8451 6885 8463 6919
rect 8404 6879 8463 6885
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8110 6808 8116 6860
rect 8168 6808 8174 6860
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8404 6848 8432 6879
rect 8570 6876 8576 6928
rect 8628 6916 8634 6928
rect 8628 6888 8984 6916
rect 8628 6876 8634 6888
rect 8352 6820 8432 6848
rect 8352 6808 8358 6820
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8956 6857 8984 6888
rect 13170 6876 13176 6928
rect 13228 6916 13234 6928
rect 13458 6919 13516 6925
rect 13458 6916 13470 6919
rect 13228 6888 13470 6916
rect 13228 6876 13234 6888
rect 13458 6885 13470 6888
rect 13504 6885 13516 6919
rect 13458 6879 13516 6885
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 9272 6820 9413 6848
rect 9272 6808 9278 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 13722 6808 13728 6860
rect 13780 6808 13786 6860
rect 8128 6780 8156 6808
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 8128 6752 9137 6780
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 8536 6684 8677 6712
rect 8536 6672 8542 6684
rect 8665 6681 8677 6684
rect 8711 6681 8723 6715
rect 8665 6675 8723 6681
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6546 6644 6552 6656
rect 6236 6616 6552 6644
rect 6236 6604 6242 6616
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 8573 6647 8631 6653
rect 8573 6613 8585 6647
rect 8619 6644 8631 6647
rect 8938 6644 8944 6656
rect 8619 6616 8944 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 10686 6604 10692 6656
rect 10744 6604 10750 6656
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 8110 6264 8116 6316
rect 8168 6304 8174 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 8168 6276 9321 6304
rect 8168 6264 8174 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9582 6264 9588 6316
rect 9640 6264 9646 6316
rect 10870 6128 10876 6180
rect 10928 6168 10934 6180
rect 10965 6171 11023 6177
rect 10965 6168 10977 6171
rect 10928 6140 10977 6168
rect 10928 6128 10934 6140
rect 10965 6137 10977 6140
rect 11011 6168 11023 6171
rect 11146 6168 11152 6180
rect 11011 6140 11152 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11146 6128 11152 6140
rect 11204 6128 11210 6180
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 13630 5556 13636 5568
rect 10744 5528 13636 5556
rect 10744 5516 10750 5528
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 1210 3340 1216 3392
rect 1268 3380 1274 3392
rect 6638 3380 6644 3392
rect 1268 3352 6644 3380
rect 1268 3340 1274 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 848 18776 900 18828
rect 2504 18776 2556 18828
rect 4160 18776 4212 18828
rect 5816 18776 5868 18828
rect 7472 18776 7524 18828
rect 9496 18844 9548 18896
rect 9128 18776 9180 18828
rect 10784 18776 10836 18828
rect 12440 18776 12492 18828
rect 14096 18776 14148 18828
rect 15752 18776 15804 18828
rect 17408 18776 17460 18828
rect 6920 18708 6972 18760
rect 6276 18640 6328 18692
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 13176 18640 13228 18692
rect 5908 18572 5960 18624
rect 6644 18572 6696 18624
rect 8576 18572 8628 18624
rect 8668 18615 8720 18624
rect 8668 18581 8677 18615
rect 8677 18581 8711 18615
rect 8711 18581 8720 18615
rect 8668 18572 8720 18581
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 10876 18572 10928 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 9496 18368 9548 18420
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 8392 18207 8444 18216
rect 8392 18173 8401 18207
rect 8401 18173 8435 18207
rect 8435 18173 8444 18207
rect 8392 18164 8444 18173
rect 8668 18207 8720 18216
rect 8668 18173 8702 18207
rect 8702 18173 8720 18207
rect 8668 18164 8720 18173
rect 11060 18207 11112 18216
rect 11060 18173 11069 18207
rect 11069 18173 11103 18207
rect 11103 18173 11112 18207
rect 11060 18164 11112 18173
rect 12992 18164 13044 18216
rect 13084 18207 13136 18216
rect 13084 18173 13093 18207
rect 13093 18173 13127 18207
rect 13127 18173 13136 18207
rect 13084 18164 13136 18173
rect 13176 18207 13228 18216
rect 13176 18173 13185 18207
rect 13185 18173 13219 18207
rect 13219 18173 13228 18207
rect 13176 18164 13228 18173
rect 17500 18164 17552 18216
rect 6000 18096 6052 18148
rect 12348 18096 12400 18148
rect 15384 18139 15436 18148
rect 15384 18105 15393 18139
rect 15393 18105 15427 18139
rect 15427 18105 15436 18139
rect 15384 18096 15436 18105
rect 7380 18071 7432 18080
rect 7380 18037 7389 18071
rect 7389 18037 7423 18071
rect 7423 18037 7432 18071
rect 7380 18028 7432 18037
rect 9220 18028 9272 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 13728 18028 13780 18080
rect 16672 18028 16724 18080
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 6000 17867 6052 17876
rect 6000 17833 6009 17867
rect 6009 17833 6043 17867
rect 6043 17833 6052 17867
rect 6000 17824 6052 17833
rect 9312 17824 9364 17876
rect 12348 17867 12400 17876
rect 12348 17833 12357 17867
rect 12357 17833 12391 17867
rect 12391 17833 12400 17867
rect 12348 17824 12400 17833
rect 12716 17824 12768 17876
rect 15384 17824 15436 17876
rect 5908 17688 5960 17740
rect 6920 17731 6972 17740
rect 6920 17697 6929 17731
rect 6929 17697 6963 17731
rect 6963 17697 6972 17731
rect 6920 17688 6972 17697
rect 7288 17688 7340 17740
rect 6552 17620 6604 17672
rect 8392 17756 8444 17808
rect 9036 17688 9088 17740
rect 9496 17756 9548 17808
rect 13176 17756 13228 17808
rect 5448 17552 5500 17604
rect 7380 17484 7432 17536
rect 8116 17484 8168 17536
rect 8484 17552 8536 17604
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13084 17688 13136 17740
rect 13360 17731 13412 17740
rect 13360 17697 13369 17731
rect 13369 17697 13403 17731
rect 13403 17697 13412 17731
rect 13360 17688 13412 17697
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 10876 17620 10928 17672
rect 9312 17552 9364 17604
rect 10508 17552 10560 17604
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 12532 17620 12584 17672
rect 8668 17484 8720 17536
rect 9220 17527 9272 17536
rect 9220 17493 9229 17527
rect 9229 17493 9263 17527
rect 9263 17493 9272 17527
rect 9220 17484 9272 17493
rect 9588 17484 9640 17536
rect 11612 17484 11664 17536
rect 12624 17484 12676 17536
rect 13636 17484 13688 17536
rect 14004 17484 14056 17536
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 7196 17323 7248 17332
rect 7196 17289 7205 17323
rect 7205 17289 7239 17323
rect 7239 17289 7248 17323
rect 7196 17280 7248 17289
rect 8944 17280 8996 17332
rect 9036 17323 9088 17332
rect 9036 17289 9045 17323
rect 9045 17289 9079 17323
rect 9079 17289 9088 17323
rect 9036 17280 9088 17289
rect 10324 17323 10376 17332
rect 10324 17289 10333 17323
rect 10333 17289 10367 17323
rect 10367 17289 10376 17323
rect 10324 17280 10376 17289
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 11704 17280 11756 17332
rect 6644 17144 6696 17196
rect 4160 17076 4212 17128
rect 5448 17076 5500 17128
rect 6552 17119 6604 17128
rect 6552 17085 6561 17119
rect 6561 17085 6595 17119
rect 6595 17085 6604 17119
rect 6552 17076 6604 17085
rect 6920 17076 6972 17128
rect 8116 17144 8168 17196
rect 8576 17144 8628 17196
rect 7288 17076 7340 17128
rect 8024 17076 8076 17128
rect 9312 17144 9364 17196
rect 12624 17212 12676 17264
rect 9496 17076 9548 17128
rect 11428 17076 11480 17128
rect 12532 17144 12584 17196
rect 11612 17119 11664 17128
rect 11612 17085 11621 17119
rect 11621 17085 11655 17119
rect 11655 17085 11664 17119
rect 11612 17076 11664 17085
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 16672 17280 16724 17332
rect 12992 17144 13044 17196
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 12164 17076 12216 17085
rect 13084 17119 13136 17128
rect 13084 17085 13093 17119
rect 13093 17085 13127 17119
rect 13127 17085 13136 17119
rect 13084 17076 13136 17085
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 14188 17076 14240 17128
rect 10324 17008 10376 17060
rect 10784 17008 10836 17060
rect 6368 16940 6420 16992
rect 9496 16940 9548 16992
rect 11336 16940 11388 16992
rect 11520 16940 11572 16992
rect 12348 16983 12400 16992
rect 12348 16949 12357 16983
rect 12357 16949 12391 16983
rect 12391 16949 12400 16983
rect 12348 16940 12400 16949
rect 12900 16940 12952 16992
rect 13912 16940 13964 16992
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 6644 16736 6696 16788
rect 6368 16643 6420 16652
rect 6368 16609 6377 16643
rect 6377 16609 6411 16643
rect 6411 16609 6420 16643
rect 6368 16600 6420 16609
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 7196 16600 7248 16652
rect 7840 16600 7892 16652
rect 8944 16736 8996 16788
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 8024 16668 8076 16720
rect 12164 16668 12216 16720
rect 7380 16532 7432 16584
rect 8668 16643 8720 16652
rect 8668 16609 8677 16643
rect 8677 16609 8711 16643
rect 8711 16609 8720 16643
rect 8668 16600 8720 16609
rect 10600 16600 10652 16652
rect 12348 16600 12400 16652
rect 13360 16600 13412 16652
rect 13912 16643 13964 16652
rect 13912 16609 13921 16643
rect 13921 16609 13955 16643
rect 13955 16609 13964 16643
rect 13912 16600 13964 16609
rect 13084 16532 13136 16584
rect 7012 16464 7064 16516
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 8852 16439 8904 16448
rect 8852 16405 8861 16439
rect 8861 16405 8895 16439
rect 8895 16405 8904 16439
rect 8852 16396 8904 16405
rect 9220 16396 9272 16448
rect 13820 16439 13872 16448
rect 13820 16405 13829 16439
rect 13829 16405 13863 16439
rect 13863 16405 13872 16439
rect 13820 16396 13872 16405
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 6644 16124 6696 16176
rect 6276 16031 6328 16040
rect 6276 15997 6285 16031
rect 6285 15997 6319 16031
rect 6319 15997 6328 16031
rect 6276 15988 6328 15997
rect 6736 15988 6788 16040
rect 6920 16192 6972 16244
rect 7932 16192 7984 16244
rect 10324 16192 10376 16244
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7380 15988 7432 16040
rect 7840 15988 7892 16040
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 9312 16056 9364 16108
rect 9220 16031 9272 16040
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 6184 15852 6236 15904
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 9036 15963 9088 15972
rect 9036 15929 9045 15963
rect 9045 15929 9079 15963
rect 9079 15929 9088 15963
rect 9036 15920 9088 15929
rect 9128 15963 9180 15972
rect 9128 15929 9137 15963
rect 9137 15929 9171 15963
rect 9171 15929 9180 15963
rect 9128 15920 9180 15929
rect 9864 16031 9916 16040
rect 9864 15997 9873 16031
rect 9873 15997 9907 16031
rect 9907 15997 9916 16031
rect 9864 15988 9916 15997
rect 7104 15852 7156 15904
rect 7380 15895 7432 15904
rect 7380 15861 7389 15895
rect 7389 15861 7423 15895
rect 7423 15861 7432 15895
rect 7380 15852 7432 15861
rect 8576 15852 8628 15904
rect 10784 15988 10836 16040
rect 11152 16124 11204 16176
rect 12624 16124 12676 16176
rect 13452 16056 13504 16108
rect 12532 15988 12584 16040
rect 13728 16031 13780 16040
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 14004 16031 14056 16040
rect 14004 15997 14013 16031
rect 14013 15997 14047 16031
rect 14047 15997 14056 16031
rect 14004 15988 14056 15997
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 10508 15852 10560 15904
rect 12440 15895 12492 15904
rect 12440 15861 12449 15895
rect 12449 15861 12483 15895
rect 12483 15861 12492 15895
rect 12440 15852 12492 15861
rect 12992 15852 13044 15904
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 6920 15648 6972 15700
rect 9036 15648 9088 15700
rect 9128 15691 9180 15700
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 5080 15512 5132 15564
rect 6368 15512 6420 15564
rect 7288 15580 7340 15632
rect 7380 15623 7432 15632
rect 7380 15589 7389 15623
rect 7389 15589 7423 15623
rect 7423 15589 7432 15623
rect 7380 15580 7432 15589
rect 8852 15623 8904 15632
rect 8852 15589 8861 15623
rect 8861 15589 8895 15623
rect 8895 15589 8904 15623
rect 8852 15580 8904 15589
rect 7012 15512 7064 15564
rect 4160 15444 4212 15496
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 7380 15444 7432 15496
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 13544 15648 13596 15700
rect 14924 15648 14976 15700
rect 12440 15580 12492 15632
rect 9588 15444 9640 15496
rect 10508 15555 10560 15564
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 11060 15512 11112 15564
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 10968 15487 11020 15496
rect 10968 15453 10977 15487
rect 10977 15453 11011 15487
rect 11011 15453 11020 15487
rect 10968 15444 11020 15453
rect 7196 15376 7248 15428
rect 10232 15376 10284 15428
rect 5632 15351 5684 15360
rect 5632 15317 5641 15351
rect 5641 15317 5675 15351
rect 5675 15317 5684 15351
rect 5632 15308 5684 15317
rect 9312 15308 9364 15360
rect 11152 15308 11204 15360
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 5080 15147 5132 15156
rect 5080 15113 5089 15147
rect 5089 15113 5123 15147
rect 5123 15113 5132 15147
rect 5080 15104 5132 15113
rect 6644 15104 6696 15156
rect 9680 15104 9732 15156
rect 11060 15104 11112 15156
rect 12256 15104 12308 15156
rect 13452 15104 13504 15156
rect 6736 15079 6788 15088
rect 6736 15045 6745 15079
rect 6745 15045 6779 15079
rect 6779 15045 6788 15079
rect 6736 15036 6788 15045
rect 6828 15036 6880 15088
rect 7196 15036 7248 15088
rect 5448 14900 5500 14952
rect 5632 14900 5684 14952
rect 6828 14900 6880 14952
rect 7840 14968 7892 15020
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 7380 14943 7432 14952
rect 7380 14909 7389 14943
rect 7389 14909 7423 14943
rect 7423 14909 7432 14943
rect 7380 14900 7432 14909
rect 8024 14900 8076 14952
rect 10416 14900 10468 14952
rect 6092 14807 6144 14816
rect 6092 14773 6101 14807
rect 6101 14773 6135 14807
rect 6135 14773 6144 14807
rect 6092 14764 6144 14773
rect 6552 14764 6604 14816
rect 8576 14832 8628 14884
rect 10784 14832 10836 14884
rect 7196 14764 7248 14816
rect 7288 14807 7340 14816
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 7380 14764 7432 14816
rect 8116 14764 8168 14816
rect 12072 14764 12124 14816
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 4160 14560 4212 14612
rect 6828 14560 6880 14612
rect 8852 14560 8904 14612
rect 5448 14356 5500 14408
rect 6552 14535 6604 14544
rect 6552 14501 6561 14535
rect 6561 14501 6595 14535
rect 6595 14501 6604 14535
rect 6552 14492 6604 14501
rect 10416 14603 10468 14612
rect 10416 14569 10425 14603
rect 10425 14569 10459 14603
rect 10459 14569 10468 14603
rect 10416 14560 10468 14569
rect 12164 14560 12216 14612
rect 12256 14603 12308 14612
rect 12256 14569 12265 14603
rect 12265 14569 12299 14603
rect 12299 14569 12308 14603
rect 12256 14560 12308 14569
rect 6184 14288 6236 14340
rect 6644 14399 6696 14408
rect 6644 14365 6653 14399
rect 6653 14365 6687 14399
rect 6687 14365 6696 14399
rect 6644 14356 6696 14365
rect 6828 14356 6880 14408
rect 8208 14356 8260 14408
rect 8760 14467 8812 14476
rect 8760 14433 8769 14467
rect 8769 14433 8803 14467
rect 8803 14433 8812 14467
rect 8760 14424 8812 14433
rect 9128 14424 9180 14476
rect 9956 14424 10008 14476
rect 10784 14535 10836 14544
rect 10784 14501 10793 14535
rect 10793 14501 10827 14535
rect 10827 14501 10836 14535
rect 10784 14492 10836 14501
rect 11704 14535 11756 14544
rect 11704 14501 11713 14535
rect 11713 14501 11747 14535
rect 11747 14501 11756 14535
rect 11704 14492 11756 14501
rect 11152 14467 11204 14476
rect 11152 14433 11161 14467
rect 11161 14433 11195 14467
rect 11195 14433 11204 14467
rect 11152 14424 11204 14433
rect 6368 14288 6420 14340
rect 9772 14356 9824 14408
rect 11060 14356 11112 14408
rect 12348 14424 12400 14476
rect 12532 14424 12584 14476
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 13084 14492 13136 14544
rect 13452 14492 13504 14544
rect 12992 14356 13044 14408
rect 12164 14288 12216 14340
rect 12440 14288 12492 14340
rect 12716 14288 12768 14340
rect 12808 14331 12860 14340
rect 12808 14297 12817 14331
rect 12817 14297 12851 14331
rect 12851 14297 12860 14331
rect 12808 14288 12860 14297
rect 6092 14220 6144 14272
rect 8116 14220 8168 14272
rect 8576 14220 8628 14272
rect 9312 14220 9364 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 11704 14220 11756 14272
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 7012 14016 7064 14068
rect 7104 14016 7156 14068
rect 6736 13948 6788 14000
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 7104 13880 7156 13932
rect 8208 13923 8260 13932
rect 8208 13889 8217 13923
rect 8217 13889 8251 13923
rect 8251 13889 8260 13923
rect 8208 13880 8260 13889
rect 4160 13812 4212 13864
rect 6184 13855 6236 13864
rect 6184 13821 6193 13855
rect 6193 13821 6227 13855
rect 6227 13821 6236 13855
rect 6184 13812 6236 13821
rect 6552 13855 6604 13864
rect 6552 13821 6561 13855
rect 6561 13821 6595 13855
rect 6595 13821 6604 13855
rect 6552 13812 6604 13821
rect 5632 13744 5684 13796
rect 8576 13855 8628 13864
rect 8576 13821 8585 13855
rect 8585 13821 8619 13855
rect 8619 13821 8628 13855
rect 8576 13812 8628 13821
rect 9128 13948 9180 14000
rect 9772 14016 9824 14068
rect 10232 14016 10284 14068
rect 12072 14016 12124 14068
rect 12440 14016 12492 14068
rect 12624 14016 12676 14068
rect 13084 14016 13136 14068
rect 11704 13948 11756 14000
rect 7288 13744 7340 13796
rect 7656 13744 7708 13796
rect 9128 13855 9180 13864
rect 9128 13821 9137 13855
rect 9137 13821 9171 13855
rect 9171 13821 9180 13855
rect 9128 13812 9180 13821
rect 9680 13880 9732 13932
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 11520 13880 11572 13932
rect 12532 13948 12584 14000
rect 12716 13948 12768 14000
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 9588 13744 9640 13796
rect 9956 13744 10008 13796
rect 8852 13676 8904 13728
rect 12164 13855 12216 13864
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 11704 13787 11756 13796
rect 11704 13753 11713 13787
rect 11713 13753 11747 13787
rect 11747 13753 11756 13787
rect 11704 13744 11756 13753
rect 11796 13744 11848 13796
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 12716 13855 12768 13864
rect 12716 13821 12725 13855
rect 12725 13821 12759 13855
rect 12759 13821 12768 13855
rect 12716 13812 12768 13821
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 12992 13855 13044 13864
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 12532 13676 12584 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 6552 13472 6604 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 8760 13515 8812 13524
rect 8760 13481 8795 13515
rect 8795 13481 8812 13515
rect 8760 13472 8812 13481
rect 9588 13472 9640 13524
rect 11152 13472 11204 13524
rect 12164 13472 12216 13524
rect 12624 13472 12676 13524
rect 12808 13472 12860 13524
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 7012 13404 7064 13456
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 7380 13336 7432 13388
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7380 13200 7432 13252
rect 8116 13200 8168 13252
rect 9680 13404 9732 13456
rect 11520 13404 11572 13456
rect 12072 13404 12124 13456
rect 10968 13336 11020 13388
rect 11704 13268 11756 13320
rect 12992 13268 13044 13320
rect 9312 13200 9364 13252
rect 12716 13200 12768 13252
rect 8852 13132 8904 13184
rect 8944 13175 8996 13184
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 6828 12928 6880 12980
rect 9128 12971 9180 12980
rect 9128 12937 9137 12971
rect 9137 12937 9171 12971
rect 9171 12937 9180 12971
rect 9128 12928 9180 12937
rect 9312 12928 9364 12980
rect 9588 12928 9640 12980
rect 11060 12928 11112 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 11796 12928 11848 12980
rect 13084 12928 13136 12980
rect 6184 12792 6236 12844
rect 4988 12631 5040 12640
rect 4988 12597 4997 12631
rect 4997 12597 5031 12631
rect 5031 12597 5040 12631
rect 4988 12588 5040 12597
rect 5540 12724 5592 12776
rect 5632 12767 5684 12776
rect 5632 12733 5641 12767
rect 5641 12733 5675 12767
rect 5675 12733 5684 12767
rect 5632 12724 5684 12733
rect 6460 12699 6512 12708
rect 6460 12665 6469 12699
rect 6469 12665 6503 12699
rect 6503 12665 6512 12699
rect 6460 12656 6512 12665
rect 6552 12588 6604 12640
rect 6644 12631 6696 12640
rect 8944 12792 8996 12844
rect 8392 12724 8444 12776
rect 8576 12724 8628 12776
rect 9588 12792 9640 12844
rect 11704 12792 11756 12844
rect 11888 12792 11940 12844
rect 10324 12724 10376 12776
rect 11152 12724 11204 12776
rect 12532 12860 12584 12912
rect 12992 12792 13044 12844
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 13084 12724 13136 12776
rect 6644 12597 6669 12631
rect 6669 12597 6696 12631
rect 6644 12588 6696 12597
rect 8852 12588 8904 12640
rect 9588 12588 9640 12640
rect 13912 12656 13964 12708
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 5540 12384 5592 12436
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 7380 12384 7432 12436
rect 7840 12384 7892 12436
rect 7932 12384 7984 12436
rect 9588 12384 9640 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 4988 12316 5040 12368
rect 6736 12316 6788 12368
rect 8760 12316 8812 12368
rect 4160 12291 4212 12300
rect 4160 12257 4169 12291
rect 4169 12257 4203 12291
rect 4203 12257 4212 12291
rect 4160 12248 4212 12257
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 6644 12248 6696 12300
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 6368 12180 6420 12232
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 7748 12291 7800 12300
rect 7748 12257 7757 12291
rect 7757 12257 7791 12291
rect 7791 12257 7800 12291
rect 7748 12248 7800 12257
rect 8116 12248 8168 12300
rect 8208 12248 8260 12300
rect 10968 12316 11020 12368
rect 12900 12384 12952 12436
rect 13084 12384 13136 12436
rect 12716 12359 12768 12368
rect 12716 12325 12725 12359
rect 12725 12325 12759 12359
rect 12759 12325 12768 12359
rect 12716 12316 12768 12325
rect 9588 12248 9640 12300
rect 8024 12180 8076 12232
rect 9864 12248 9916 12300
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 12072 12248 12124 12300
rect 13084 12291 13136 12300
rect 13084 12257 13093 12291
rect 13093 12257 13127 12291
rect 13127 12257 13136 12291
rect 13084 12248 13136 12257
rect 7932 12112 7984 12164
rect 7380 12044 7432 12096
rect 7748 12044 7800 12096
rect 8208 12044 8260 12096
rect 9036 12044 9088 12096
rect 9956 12180 10008 12232
rect 10140 12112 10192 12164
rect 11152 12112 11204 12164
rect 12532 12112 12584 12164
rect 10876 12044 10928 12096
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 5908 11840 5960 11892
rect 8024 11883 8076 11892
rect 8024 11849 8033 11883
rect 8033 11849 8067 11883
rect 8067 11849 8076 11883
rect 8024 11840 8076 11849
rect 8116 11883 8168 11892
rect 8116 11849 8125 11883
rect 8125 11849 8159 11883
rect 8159 11849 8168 11883
rect 8116 11840 8168 11849
rect 8852 11840 8904 11892
rect 13636 11840 13688 11892
rect 4160 11636 4212 11688
rect 5724 11568 5776 11620
rect 6552 11704 6604 11756
rect 6460 11636 6512 11688
rect 7840 11704 7892 11756
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 6644 11568 6696 11620
rect 7472 11679 7524 11688
rect 7472 11645 7481 11679
rect 7481 11645 7515 11679
rect 7515 11645 7524 11679
rect 7472 11636 7524 11645
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 9956 11704 10008 11756
rect 12072 11772 12124 11824
rect 7932 11568 7984 11620
rect 10232 11636 10284 11688
rect 11612 11636 11664 11688
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 15108 11704 15160 11756
rect 9864 11568 9916 11620
rect 10784 11568 10836 11620
rect 11704 11568 11756 11620
rect 6092 11500 6144 11552
rect 6276 11500 6328 11552
rect 6736 11500 6788 11552
rect 7472 11500 7524 11552
rect 8760 11543 8812 11552
rect 8760 11509 8769 11543
rect 8769 11509 8803 11543
rect 8803 11509 8812 11543
rect 8760 11500 8812 11509
rect 9680 11500 9732 11552
rect 10324 11500 10376 11552
rect 10968 11500 11020 11552
rect 11152 11500 11204 11552
rect 11520 11500 11572 11552
rect 12992 11636 13044 11688
rect 14004 11568 14056 11620
rect 13912 11543 13964 11552
rect 13912 11509 13921 11543
rect 13921 11509 13955 11543
rect 13955 11509 13964 11543
rect 13912 11500 13964 11509
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 5724 11296 5776 11348
rect 6460 11296 6512 11348
rect 8392 11296 8444 11348
rect 9312 11296 9364 11348
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 12164 11296 12216 11348
rect 12992 11339 13044 11348
rect 12992 11305 13001 11339
rect 13001 11305 13035 11339
rect 13035 11305 13044 11339
rect 12992 11296 13044 11305
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 6368 11228 6420 11280
rect 6736 11228 6788 11280
rect 7380 11228 7432 11280
rect 10600 11228 10652 11280
rect 10968 11228 11020 11280
rect 6276 11203 6328 11212
rect 6276 11169 6285 11203
rect 6285 11169 6319 11203
rect 6319 11169 6328 11203
rect 6276 11160 6328 11169
rect 6644 11160 6696 11212
rect 11060 11160 11112 11212
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 11612 11160 11664 11212
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 12900 11228 12952 11280
rect 4160 11092 4212 11144
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 8300 11092 8352 11144
rect 8760 11135 8812 11144
rect 8760 11101 8769 11135
rect 8769 11101 8803 11135
rect 8803 11101 8812 11135
rect 8760 11092 8812 11101
rect 10232 11092 10284 11144
rect 10876 11092 10928 11144
rect 5632 11024 5684 11076
rect 6644 11024 6696 11076
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 13820 10956 13872 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 7104 10684 7156 10736
rect 6828 10548 6880 10600
rect 8208 10616 8260 10668
rect 10324 10616 10376 10668
rect 11060 10616 11112 10668
rect 7932 10591 7984 10600
rect 7932 10557 7941 10591
rect 7941 10557 7975 10591
rect 7975 10557 7984 10591
rect 7932 10548 7984 10557
rect 10232 10548 10284 10600
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 6184 10412 6236 10464
rect 6552 10412 6604 10464
rect 6736 10412 6788 10464
rect 7840 10480 7892 10532
rect 12624 10548 12676 10600
rect 14004 10616 14056 10668
rect 11888 10480 11940 10532
rect 11704 10455 11756 10464
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 15660 10548 15712 10600
rect 13820 10412 13872 10464
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 18604 10412 18656 10464
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 5540 10140 5592 10192
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 6828 10208 6880 10260
rect 6736 10115 6788 10124
rect 4988 9868 5040 9920
rect 5816 9868 5868 9920
rect 6184 9868 6236 9920
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7380 10140 7432 10192
rect 9220 10183 9272 10192
rect 9220 10149 9229 10183
rect 9229 10149 9263 10183
rect 9263 10149 9272 10183
rect 9220 10140 9272 10149
rect 9496 10208 9548 10260
rect 12624 10208 12676 10260
rect 12716 10251 12768 10260
rect 12716 10217 12725 10251
rect 12725 10217 12759 10251
rect 12759 10217 12768 10251
rect 12716 10208 12768 10217
rect 12808 10208 12860 10260
rect 12532 10140 12584 10192
rect 7932 10072 7984 10124
rect 10232 10072 10284 10124
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10416 10072 10468 10124
rect 7840 10004 7892 10056
rect 12716 10072 12768 10124
rect 13912 10072 13964 10124
rect 13084 10004 13136 10056
rect 13820 10004 13872 10056
rect 7288 9979 7340 9988
rect 7288 9945 7297 9979
rect 7297 9945 7331 9979
rect 7331 9945 7340 9979
rect 7288 9936 7340 9945
rect 8024 9936 8076 9988
rect 10508 9936 10560 9988
rect 12992 9979 13044 9988
rect 12992 9945 13001 9979
rect 13001 9945 13035 9979
rect 13035 9945 13044 9979
rect 12992 9936 13044 9945
rect 6368 9868 6420 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 8944 9868 8996 9920
rect 9772 9868 9824 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11244 9868 11296 9920
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 13268 9868 13320 9877
rect 14096 9868 14148 9920
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 16120 9868 16172 9920
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 6092 9664 6144 9716
rect 9220 9664 9272 9716
rect 10416 9707 10468 9716
rect 10416 9673 10425 9707
rect 10425 9673 10459 9707
rect 10459 9673 10468 9707
rect 10416 9664 10468 9673
rect 10692 9664 10744 9716
rect 6184 9596 6236 9648
rect 4160 9528 4212 9580
rect 8944 9571 8996 9580
rect 8944 9537 8953 9571
rect 8953 9537 8987 9571
rect 8987 9537 8996 9571
rect 8944 9528 8996 9537
rect 9772 9596 9824 9648
rect 12808 9639 12860 9648
rect 12808 9605 12817 9639
rect 12817 9605 12851 9639
rect 12851 9605 12860 9639
rect 12808 9596 12860 9605
rect 6184 9460 6236 9512
rect 7380 9460 7432 9512
rect 9128 9528 9180 9580
rect 4896 9392 4948 9444
rect 7196 9392 7248 9444
rect 7472 9392 7524 9444
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 9588 9528 9640 9580
rect 10232 9528 10284 9580
rect 10600 9528 10652 9580
rect 11888 9528 11940 9580
rect 12164 9571 12216 9580
rect 12164 9537 12173 9571
rect 12173 9537 12207 9571
rect 12207 9537 12216 9571
rect 12164 9528 12216 9537
rect 12348 9528 12400 9580
rect 12716 9528 12768 9580
rect 9864 9392 9916 9444
rect 10416 9460 10468 9512
rect 10692 9503 10744 9512
rect 10692 9469 10701 9503
rect 10701 9469 10735 9503
rect 10735 9469 10744 9503
rect 10692 9460 10744 9469
rect 10876 9392 10928 9444
rect 12440 9460 12492 9512
rect 12532 9503 12584 9512
rect 12532 9469 12541 9503
rect 12541 9469 12575 9503
rect 12575 9469 12584 9503
rect 12532 9460 12584 9469
rect 13084 9460 13136 9512
rect 12992 9392 13044 9444
rect 13360 9503 13412 9512
rect 13360 9469 13369 9503
rect 13369 9469 13403 9503
rect 13403 9469 13412 9503
rect 13360 9460 13412 9469
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 6460 9324 6512 9376
rect 8392 9324 8444 9376
rect 8852 9367 8904 9376
rect 8852 9333 8861 9367
rect 8861 9333 8895 9367
rect 8895 9333 8904 9367
rect 8852 9324 8904 9333
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 9404 9324 9456 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10324 9324 10376 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 11888 9367 11940 9376
rect 11888 9333 11913 9367
rect 11913 9333 11940 9367
rect 11888 9324 11940 9333
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 12900 9324 12952 9376
rect 13820 9392 13872 9444
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 4896 9120 4948 9172
rect 5540 9120 5592 9172
rect 7472 9120 7524 9172
rect 9220 9120 9272 9172
rect 10692 9120 10744 9172
rect 11888 9120 11940 9172
rect 13268 9120 13320 9172
rect 13820 9120 13872 9172
rect 6092 9052 6144 9104
rect 6552 9095 6604 9104
rect 6552 9061 6561 9095
rect 6561 9061 6595 9095
rect 6595 9061 6604 9095
rect 6552 9052 6604 9061
rect 4988 8984 5040 9036
rect 6368 8984 6420 9036
rect 6736 8984 6788 9036
rect 6920 9052 6972 9104
rect 8852 9052 8904 9104
rect 6460 8916 6512 8968
rect 7104 8984 7156 9036
rect 7196 9027 7248 9036
rect 7196 8993 7205 9027
rect 7205 8993 7239 9027
rect 7239 8993 7248 9027
rect 7196 8984 7248 8993
rect 8024 8984 8076 9036
rect 9128 8984 9180 9036
rect 9312 8984 9364 9036
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 10508 9052 10560 9104
rect 12072 9052 12124 9104
rect 14096 9095 14148 9104
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10232 8984 10284 9036
rect 12624 8984 12676 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 13084 9027 13136 9036
rect 12716 8984 12768 8993
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 13360 8984 13412 9036
rect 14096 9061 14130 9095
rect 14130 9061 14148 9095
rect 14096 9052 14148 9061
rect 6276 8848 6328 8900
rect 6828 8848 6880 8900
rect 8392 8916 8444 8968
rect 11152 8916 11204 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12164 8848 12216 8900
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 9220 8823 9272 8832
rect 9220 8789 9229 8823
rect 9229 8789 9263 8823
rect 9263 8789 9272 8823
rect 9220 8780 9272 8789
rect 13084 8848 13136 8900
rect 13728 8916 13780 8968
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 6092 8372 6144 8424
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 6276 8415 6328 8424
rect 6276 8381 6285 8415
rect 6285 8381 6319 8415
rect 6319 8381 6328 8415
rect 6276 8372 6328 8381
rect 7656 8576 7708 8628
rect 9496 8576 9548 8628
rect 9680 8576 9732 8628
rect 9864 8576 9916 8628
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 12900 8576 12952 8628
rect 13084 8576 13136 8628
rect 10784 8508 10836 8560
rect 12624 8508 12676 8560
rect 9312 8440 9364 8492
rect 6644 8372 6696 8424
rect 7288 8372 7340 8424
rect 8760 8415 8812 8424
rect 8760 8381 8769 8415
rect 8769 8381 8803 8415
rect 8803 8381 8812 8415
rect 8760 8372 8812 8381
rect 8944 8415 8996 8424
rect 8944 8381 8953 8415
rect 8953 8381 8987 8415
rect 8987 8381 8996 8415
rect 8944 8372 8996 8381
rect 9128 8372 9180 8424
rect 10692 8372 10744 8424
rect 11060 8415 11112 8424
rect 11060 8381 11069 8415
rect 11069 8381 11103 8415
rect 11103 8381 11112 8415
rect 11060 8372 11112 8381
rect 8300 8304 8352 8356
rect 6276 8236 6328 8288
rect 6736 8236 6788 8288
rect 9312 8304 9364 8356
rect 12716 8347 12768 8356
rect 12716 8313 12725 8347
rect 12725 8313 12759 8347
rect 12759 8313 12768 8347
rect 12716 8304 12768 8313
rect 9128 8236 9180 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 13360 8236 13412 8288
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 11060 8032 11112 8084
rect 11336 8032 11388 8084
rect 12072 8032 12124 8084
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8024 7871 8076 7880
rect 8024 7837 8033 7871
rect 8033 7837 8067 7871
rect 8067 7837 8076 7871
rect 8024 7828 8076 7837
rect 8208 7896 8260 7948
rect 8576 7828 8628 7880
rect 8760 7939 8812 7948
rect 8760 7905 8769 7939
rect 8769 7905 8803 7939
rect 8803 7905 8812 7939
rect 8760 7896 8812 7905
rect 9036 7939 9088 7948
rect 9036 7905 9045 7939
rect 9045 7905 9079 7939
rect 9079 7905 9088 7939
rect 9036 7896 9088 7905
rect 9128 7939 9180 7948
rect 9128 7905 9137 7939
rect 9137 7905 9171 7939
rect 9171 7905 9180 7939
rect 9128 7896 9180 7905
rect 9312 7939 9364 7948
rect 9312 7905 9321 7939
rect 9321 7905 9355 7939
rect 9355 7905 9364 7939
rect 9312 7896 9364 7905
rect 10232 7964 10284 8016
rect 12532 8007 12584 8016
rect 9496 7896 9548 7948
rect 8852 7828 8904 7880
rect 10784 7896 10836 7948
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 12532 7973 12541 8007
rect 12541 7973 12575 8007
rect 12575 7973 12584 8007
rect 12532 7964 12584 7973
rect 11244 7828 11296 7880
rect 12808 7896 12860 7948
rect 13176 7896 13228 7948
rect 6276 7692 6328 7744
rect 7840 7692 7892 7744
rect 8484 7692 8536 7744
rect 8668 7692 8720 7744
rect 8944 7692 8996 7744
rect 9496 7692 9548 7744
rect 10968 7760 11020 7812
rect 12624 7692 12676 7744
rect 12716 7735 12768 7744
rect 12716 7701 12725 7735
rect 12725 7701 12759 7735
rect 12759 7701 12768 7735
rect 12716 7692 12768 7701
rect 12900 7692 12952 7744
rect 13360 7828 13412 7880
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 6552 7488 6604 7540
rect 6828 7488 6880 7540
rect 8576 7488 8628 7540
rect 10968 7531 11020 7540
rect 10968 7497 10977 7531
rect 10977 7497 11011 7531
rect 11011 7497 11020 7531
rect 10968 7488 11020 7497
rect 6276 7395 6328 7404
rect 6276 7361 6285 7395
rect 6285 7361 6319 7395
rect 6319 7361 6328 7395
rect 6276 7352 6328 7361
rect 7380 7352 7432 7404
rect 8116 7352 8168 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 8852 7352 8904 7404
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 6828 7284 6880 7336
rect 3700 7216 3752 7268
rect 6552 7216 6604 7268
rect 7104 7148 7156 7200
rect 8392 7216 8444 7268
rect 8668 7148 8720 7200
rect 8760 7148 8812 7200
rect 13728 7352 13780 7404
rect 11152 7284 11204 7336
rect 11704 7216 11756 7268
rect 12624 7327 12676 7336
rect 12624 7293 12633 7327
rect 12633 7293 12667 7327
rect 12667 7293 12676 7327
rect 12624 7284 12676 7293
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 12900 7284 12952 7336
rect 12532 7216 12584 7268
rect 12808 7148 12860 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 6552 6944 6604 6996
rect 9680 6944 9732 6996
rect 12532 6944 12584 6996
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 8300 6808 8352 6860
rect 8576 6876 8628 6928
rect 8668 6851 8720 6860
rect 8668 6817 8677 6851
rect 8677 6817 8711 6851
rect 8711 6817 8720 6851
rect 8668 6808 8720 6817
rect 13176 6876 13228 6928
rect 9220 6808 9272 6860
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 8484 6672 8536 6724
rect 6184 6604 6236 6656
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8944 6604 8996 6656
rect 10692 6647 10744 6656
rect 10692 6613 10701 6647
rect 10701 6613 10735 6647
rect 10735 6613 10744 6647
rect 10692 6604 10744 6613
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 8116 6264 8168 6316
rect 9588 6307 9640 6316
rect 9588 6273 9597 6307
rect 9597 6273 9631 6307
rect 9631 6273 9640 6307
rect 9588 6264 9640 6273
rect 10876 6128 10928 6180
rect 11152 6128 11204 6180
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 10692 5516 10744 5568
rect 13636 5516 13688 5568
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 1216 3340 1268 3392
rect 6644 3340 6696 3392
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 846 19600 902 20000
rect 2502 19600 2558 20000
rect 4158 19600 4214 20000
rect 5814 19600 5870 20000
rect 7470 19600 7526 20000
rect 9126 19600 9182 20000
rect 10782 19600 10838 20000
rect 12438 19600 12494 20000
rect 14094 19600 14150 20000
rect 15750 19600 15806 20000
rect 17406 19600 17462 20000
rect 19062 19600 19118 20000
rect 860 18834 888 19600
rect 2516 18834 2544 19600
rect 4172 18834 4200 19600
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 5828 18834 5856 19600
rect 7484 18834 7512 19600
rect 9140 18834 9168 19600
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 9496 18896 9548 18902
rect 9496 18838 9548 18844
rect 848 18828 900 18834
rect 848 18770 900 18776
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 2755 18459 3063 18468
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 5460 17610 5488 18158
rect 5920 17746 5948 18566
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6012 17882 6040 18090
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 5460 17134 5488 17546
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 4172 15502 4200 17070
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 4172 14618 4200 15438
rect 5092 15162 5120 15506
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5080 15156 5132 15162
rect 5080 15098 5132 15104
rect 5644 14958 5672 15302
rect 5448 14952 5500 14958
rect 5448 14894 5500 14900
rect 5632 14952 5684 14958
rect 5632 14894 5684 14900
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 4172 13870 4200 14554
rect 5460 14414 5488 14894
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 4172 12306 4200 13806
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 5644 12782 5672 13738
rect 5540 12776 5592 12782
rect 5540 12718 5592 12724
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 12374 5028 12582
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 5552 12442 5580 12718
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4172 11150 4200 11630
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 4172 9586 4200 11086
rect 5644 11082 5672 12718
rect 5920 11898 5948 17682
rect 6288 16046 6316 18634
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 17134 6592 17614
rect 6656 17202 6684 18566
rect 6932 18222 6960 18702
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 6932 17746 6960 18158
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6380 16658 6408 16934
rect 6656 16794 6684 17138
rect 6932 17134 6960 17682
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 7208 16658 7236 17274
rect 7300 17134 7328 17682
rect 7392 17542 7420 18022
rect 8404 17814 8432 18158
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14278 6132 14758
rect 6196 14346 6224 15846
rect 6380 15570 6408 16594
rect 6932 16250 6960 16594
rect 7300 16538 7328 17070
rect 7392 16590 7420 17478
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 8128 17202 8156 17478
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16726 8064 17070
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 7116 16510 7328 16538
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6656 15162 6684 16118
rect 7024 16046 7052 16458
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14550 6592 14758
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6656 14414 6684 15098
rect 6748 15094 6776 15982
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15706 6960 15914
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 7024 15570 7052 15982
rect 7116 15910 7144 16510
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6368 14340 6420 14346
rect 6368 14282 6420 14288
rect 6092 14272 6144 14278
rect 6092 14214 6144 14220
rect 6380 13938 6408 14282
rect 6748 14006 6776 15030
rect 6840 14958 6868 15030
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6840 14414 6868 14554
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 7024 14074 7052 15506
rect 7208 15434 7236 16390
rect 7392 16046 7420 16526
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 7852 16046 7880 16594
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 16046 7972 16186
rect 7380 16040 7432 16046
rect 7300 16000 7380 16028
rect 7300 15638 7328 16000
rect 7380 15982 7432 15988
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7392 15638 7420 15846
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7380 15496 7432 15502
rect 7380 15438 7432 15444
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 7208 14822 7236 15030
rect 7392 14958 7420 15438
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6196 13394 6224 13806
rect 6564 13530 6592 13806
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 7024 13462 7052 14010
rect 7116 13938 7144 14010
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7116 13394 7144 13874
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6196 12306 6224 12786
rect 6380 12434 6408 13262
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6288 12406 6408 12434
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5908 11892 5960 11898
rect 5908 11834 5960 11840
rect 6288 11642 6316 12406
rect 6472 12238 6500 12650
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6380 11778 6408 12174
rect 6380 11750 6500 11778
rect 6564 11762 6592 12582
rect 6656 12434 6684 12582
rect 6656 12406 6776 12434
rect 6748 12374 6776 12406
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6472 11694 6500 11750
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 6196 11614 6316 11642
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 5736 11354 5764 11562
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 6104 11218 6132 11494
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 6196 10470 6224 11614
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11218 6316 11494
rect 6472 11354 6500 11630
rect 6656 11626 6684 12242
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6748 11558 6776 12310
rect 6840 12306 6868 12922
rect 7208 12442 7236 14758
rect 7300 13802 7328 14758
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7300 13326 7328 13738
rect 7392 13394 7420 14758
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13530 7696 13738
rect 7852 13530 7880 14962
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7380 13252 7432 13258
rect 7380 13194 7432 13200
rect 7392 12442 7420 13194
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 7944 12442 7972 13330
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7932 12436 7984 12442
rect 8036 12434 8064 14894
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14278 8156 14758
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 13258 8156 14214
rect 8220 13938 8248 14350
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8036 12406 8248 12434
rect 7932 12378 7984 12384
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7760 12102 7788 12242
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6748 11286 6776 11494
rect 7392 11286 7420 12038
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 7852 11762 7880 12378
rect 7944 12170 7972 12378
rect 8220 12306 8248 12406
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7484 11558 7512 11630
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 6276 11212 6328 11218
rect 6276 11154 6328 11160
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 4988 9920 5040 9926
rect 4988 9862 5040 9868
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 4908 9178 4936 9386
rect 4896 9172 4948 9178
rect 4896 9114 4948 9120
rect 5000 9042 5028 9862
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 5552 9178 5580 10134
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 5828 8634 5856 9862
rect 6104 9722 6132 10134
rect 6380 9926 6408 11222
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 11082 6684 11154
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10062 6592 10406
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6104 9110 6132 9658
rect 6196 9654 6224 9862
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6196 9518 6224 9590
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 6104 8430 6132 9046
rect 6196 8430 6224 9454
rect 6380 9042 6408 9862
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6472 8974 6500 9318
rect 6564 9110 6592 9998
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6288 8430 6316 8842
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 6288 7954 6316 8230
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 6288 7410 6316 7686
rect 6564 7546 6592 9046
rect 6656 9024 6684 11018
rect 7104 10736 7156 10742
rect 7104 10678 7156 10684
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6748 10130 6776 10406
rect 6840 10266 6868 10542
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6736 9036 6788 9042
rect 6656 8996 6736 9024
rect 6736 8978 6788 8984
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6656 7342 6684 8366
rect 6748 8294 6776 8978
rect 6840 8906 6868 10202
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9110 6960 9862
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 7116 9042 7144 10678
rect 7392 10198 7420 11086
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 7852 10538 7880 11698
rect 7944 11626 7972 12106
rect 8036 11898 8064 12174
rect 8128 11898 8156 12242
rect 8220 12102 8248 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 11694 8248 12038
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 7932 11620 7984 11626
rect 7932 11562 7984 11568
rect 7944 10962 7972 11562
rect 7944 10934 8064 10962
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9042 7236 9386
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 7300 8430 7328 9930
rect 7392 9518 7420 10134
rect 7852 10062 7880 10474
rect 7944 10130 7972 10542
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 8036 9994 8064 10934
rect 8220 10674 8248 11630
rect 8404 11354 8432 12718
rect 8496 12434 8524 17546
rect 8588 17202 8616 18566
rect 8680 18222 8708 18566
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8680 16658 8708 17478
rect 9048 17338 9076 17682
rect 9232 17542 9260 18022
rect 9324 17882 9352 18702
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8956 16794 8984 17274
rect 9324 17202 9352 17546
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8588 15570 8616 15846
rect 8864 15638 8892 16390
rect 8852 15632 8904 15638
rect 8852 15574 8904 15580
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 14890 8616 15506
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8588 14278 8616 14826
rect 8864 14618 8892 15574
rect 8956 15570 8984 16730
rect 9220 16448 9272 16454
rect 9220 16390 9272 16396
rect 9232 16046 9260 16390
rect 9312 16108 9364 16114
rect 9312 16050 9364 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 9036 15972 9088 15978
rect 9036 15914 9088 15920
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9048 15706 9076 15914
rect 9140 15706 9168 15914
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9324 15366 9352 16050
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8576 13864 8628 13870
rect 8772 13841 8800 14418
rect 9140 14006 9168 14418
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9324 13870 9352 14214
rect 9128 13864 9180 13870
rect 8576 13806 8628 13812
rect 8758 13832 8814 13841
rect 8588 12782 8616 13806
rect 9128 13806 9180 13812
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 8758 13767 8814 13776
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8496 12406 8708 12434
rect 8680 12186 8708 12406
rect 8772 12374 8800 13466
rect 8864 13190 8892 13670
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8864 12646 8892 13126
rect 8956 12850 8984 13126
rect 9140 12986 9168 13806
rect 9324 13258 9352 13806
rect 9312 13252 9364 13258
rect 9312 13194 9364 13200
rect 9324 12986 9352 13194
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8680 12158 9168 12186
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8864 11762 8892 11834
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8772 11150 8800 11494
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 7342 6868 7482
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 3700 7268 3752 7274
rect 3700 7210 3752 7216
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 1216 3392 1268 3398
rect 1216 3334 1268 3340
rect 1228 400 1256 3334
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 3712 400 3740 7210
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 6564 7002 6592 7210
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6564 6662 6592 6938
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 6196 400 6224 6598
rect 6656 3398 6684 7278
rect 7116 7206 7144 7822
rect 7392 7410 7420 9454
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7484 9178 7512 9386
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7668 7886 7696 8570
rect 8036 7886 8064 8978
rect 8220 7954 8248 10610
rect 8312 8362 8340 11086
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8956 9586 8984 9862
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8404 8974 8432 9318
rect 8864 9110 8892 9318
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7852 6866 7880 7686
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 6866 8156 7346
rect 8312 6866 8340 8298
rect 8772 7954 8800 8366
rect 8760 7948 8812 7954
rect 8760 7890 8812 7896
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 8128 6322 8156 6802
rect 8404 6662 8432 7210
rect 8496 6730 8524 7686
rect 8588 7546 8616 7822
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8588 6934 8616 7482
rect 8680 7410 8708 7686
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8772 7206 8800 7890
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 7410 8892 7822
rect 8956 7750 8984 8366
rect 9048 7954 9076 12038
rect 9140 9586 9168 12158
rect 9416 11694 9444 18566
rect 9508 18426 9536 18838
rect 10796 18834 10824 19600
rect 12452 18834 12480 19600
rect 14108 18834 14136 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 15764 18834 15792 19600
rect 17420 18834 17448 19600
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 13176 18692 13228 18698
rect 13176 18634 13228 18640
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9508 17814 9536 18362
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 9496 17808 9548 17814
rect 9496 17750 9548 17756
rect 9508 17134 9536 17750
rect 10888 17678 10916 18566
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 11060 18216 11112 18222
rect 10980 18164 11060 18170
rect 10980 18158 11112 18164
rect 10980 18142 11100 18158
rect 12348 18148 12400 18154
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9218 10296 9274 10305
rect 9218 10231 9274 10240
rect 9232 10198 9260 10231
rect 9220 10192 9272 10198
rect 9220 10134 9272 10140
rect 9220 9716 9272 9722
rect 9220 9658 9272 9664
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9140 9042 9168 9522
rect 9232 9382 9260 9658
rect 9324 9518 9352 11290
rect 9508 10266 9536 16934
rect 9600 16028 9628 17478
rect 10520 17338 10548 17546
rect 10324 17332 10376 17338
rect 10324 17274 10376 17280
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10336 17066 10364 17274
rect 10324 17060 10376 17066
rect 10324 17002 10376 17008
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 9864 16040 9916 16046
rect 9600 16000 9864 16028
rect 9600 15502 9628 16000
rect 9864 15982 9916 15988
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 10244 15434 10272 15846
rect 10232 15428 10284 15434
rect 10232 15370 10284 15376
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9692 14498 9720 15098
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 9692 14470 9812 14498
rect 9784 14414 9812 14470
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14074 9812 14350
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9600 13530 9628 13738
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9692 13462 9720 13874
rect 9968 13802 9996 14418
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9600 12850 9628 12922
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 12442 9628 12582
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 9600 12306 9628 12378
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 11762 9904 12242
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9968 11762 9996 12174
rect 10152 12170 10180 12378
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9968 11642 9996 11698
rect 10244 11694 10272 14010
rect 10336 12782 10364 16186
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15570 10548 15846
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10428 14618 10456 14894
rect 10416 14612 10468 14618
rect 10416 14554 10468 14560
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 10336 12306 10364 12718
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 9876 11626 9996 11642
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9864 11620 9996 11626
rect 9916 11614 9996 11620
rect 9864 11562 9916 11568
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9692 10010 9720 11494
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 10244 11150 10272 11630
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10244 10606 10272 11086
rect 10336 10674 10364 11494
rect 10612 11286 10640 16594
rect 10796 16046 10824 17002
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10796 14550 10824 14826
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10888 12102 10916 17614
rect 10980 15502 11008 18142
rect 12348 18090 12400 18096
rect 12360 17882 12388 18090
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12452 17746 12480 18022
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12544 17678 12572 18566
rect 13188 18222 13216 18634
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17882 12756 18022
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 12532 17672 12584 17678
rect 12532 17614 12584 17620
rect 11612 17536 11664 17542
rect 11612 17478 11664 17484
rect 11624 17134 11652 17478
rect 11716 17338 11744 17614
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 12544 17202 12572 17614
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17270 12664 17478
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 11428 17128 11480 17134
rect 11612 17128 11664 17134
rect 11480 17076 11560 17082
rect 11428 17070 11560 17076
rect 11612 17070 11664 17076
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 11440 17054 11560 17070
rect 11532 16998 11560 17054
rect 11336 16992 11388 16998
rect 11336 16934 11388 16940
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10980 13394 11008 15438
rect 11072 15162 11100 15506
rect 11164 15366 11192 16118
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11164 14482 11192 15302
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14408 11112 14414
rect 11112 14356 11192 14362
rect 11060 14350 11192 14356
rect 11072 14334 11192 14350
rect 11164 13530 11192 14334
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11072 12434 11100 12922
rect 11164 12782 11192 13466
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10980 12406 11100 12434
rect 10980 12374 11008 12406
rect 10968 12368 11020 12374
rect 10968 12310 11020 12316
rect 11058 12336 11114 12345
rect 11058 12271 11060 12280
rect 11112 12271 11114 12280
rect 11060 12242 11112 12248
rect 11164 12170 11192 12718
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10796 11354 10824 11562
rect 11164 11558 11192 12106
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10980 11286 11008 11494
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10810 10916 11086
rect 11072 10810 11100 11154
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 10232 10600 10284 10606
rect 10692 10600 10744 10606
rect 10284 10548 10364 10554
rect 10232 10542 10364 10548
rect 10692 10542 10744 10548
rect 10244 10526 10364 10542
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 10336 10130 10364 10526
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 9692 9982 9904 10010
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9654 9812 9862
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9312 9512 9364 9518
rect 9364 9472 9536 9500
rect 9312 9454 9364 9460
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9232 9178 9260 9318
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9232 8922 9260 9114
rect 9416 9042 9444 9318
rect 9312 9036 9364 9042
rect 9312 8978 9364 8984
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9140 8894 9260 8922
rect 9140 8430 9168 8894
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 7954 9168 8230
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8680 6866 8708 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 8772 2774 8800 7142
rect 8956 6662 8984 7686
rect 9232 6866 9260 8774
rect 9324 8498 9352 8978
rect 9508 8634 9536 9472
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9324 7954 9352 8298
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7750 9536 7890
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 9600 6322 9628 9522
rect 9876 9450 9904 9982
rect 10244 9586 10272 10066
rect 10428 9722 10456 10066
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10428 9518 10456 9658
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9376 9824 9382
rect 9692 9336 9772 9364
rect 9692 9042 9720 9336
rect 10324 9376 10376 9382
rect 9772 9318 9824 9324
rect 10244 9336 10324 9364
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 10244 9042 10272 9336
rect 10324 9318 10376 9324
rect 10520 9110 10548 9930
rect 10704 9722 10732 10542
rect 11072 9926 11100 10610
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10612 9058 10640 9522
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10704 9178 10732 9454
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 10232 9036 10284 9042
rect 10612 9030 10732 9058
rect 10232 8978 10284 8984
rect 9876 8634 9904 8978
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9692 7002 9720 8570
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10244 8022 10272 8978
rect 10704 8430 10732 9030
rect 10796 8566 10824 9318
rect 10784 8560 10836 8566
rect 10784 8502 10836 8508
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10232 8016 10284 8022
rect 10232 7958 10284 7964
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 10704 6662 10732 8366
rect 10796 7954 10824 8502
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 10704 5574 10732 6598
rect 10888 6186 10916 9386
rect 11164 8974 11192 11494
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 8090 11100 8366
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7546 11008 7754
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11164 7342 11192 8230
rect 11256 7886 11284 9862
rect 11348 8090 11376 16934
rect 12176 16726 12204 17070
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12360 16658 12388 16934
rect 12348 16652 12400 16658
rect 12348 16594 12400 16600
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 12636 16182 12664 17206
rect 13004 17202 13032 18158
rect 13096 17746 13124 18158
rect 13188 17814 13216 18158
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13740 17746 13768 18022
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13096 17134 13124 17682
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 12912 16794 12940 16934
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13096 16590 13124 17070
rect 13084 16584 13136 16590
rect 13084 16526 13136 16532
rect 12624 16176 12676 16182
rect 12624 16118 12676 16124
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12452 15638 12480 15846
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11716 14278 11744 14486
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11532 13938 11560 14214
rect 12084 14074 12112 14758
rect 12268 14618 12296 15098
rect 12544 14634 12572 15982
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12452 14606 12572 14634
rect 12176 14346 12204 14554
rect 12452 14498 12480 14606
rect 12360 14482 12480 14498
rect 12636 14482 12756 14498
rect 12348 14476 12480 14482
rect 12400 14470 12480 14476
rect 12348 14418 12400 14424
rect 12452 14346 12480 14470
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12636 14476 12768 14482
rect 12636 14470 12716 14476
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 11704 14000 11756 14006
rect 11756 13960 11836 13988
rect 11704 13942 11756 13948
rect 11520 13932 11572 13938
rect 11520 13874 11572 13880
rect 11808 13802 11836 13960
rect 12164 13864 12216 13870
rect 12452 13852 12480 14010
rect 12544 14006 12572 14418
rect 12636 14074 12664 14470
rect 12716 14418 12768 14424
rect 12716 14340 12768 14346
rect 12716 14282 12768 14288
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12728 14006 12756 14282
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12820 13938 12848 14282
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12624 13864 12676 13870
rect 12452 13824 12572 13852
rect 12164 13806 12216 13812
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11520 13456 11572 13462
rect 11520 13398 11572 13404
rect 11532 12986 11560 13398
rect 11716 13326 11744 13738
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11716 12850 11744 13262
rect 11808 12986 11836 13738
rect 12176 13530 12204 13806
rect 12544 13734 12572 13824
rect 12624 13806 12676 13812
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11808 12434 11836 12922
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11716 12406 11836 12434
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11218 11560 11494
rect 11624 11218 11652 11630
rect 11716 11626 11744 12406
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11716 10470 11744 11562
rect 11900 10538 11928 12786
rect 12084 12306 12112 13398
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12544 12918 12572 13670
rect 12636 13530 12664 13806
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12728 13258 12756 13806
rect 12820 13530 12848 13874
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12072 12300 12124 12306
rect 12072 12242 12124 12248
rect 12084 11830 12112 12242
rect 12544 12170 12572 12718
rect 12912 12442 12940 15506
rect 13004 14414 13032 15846
rect 13084 14544 13136 14550
rect 13084 14486 13136 14492
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14278 13032 14350
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 13954 13032 14214
rect 13096 14074 13124 14486
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13004 13926 13124 13954
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13004 13530 13032 13806
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 13004 13326 13032 13466
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13096 12986 13124 13926
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12716 12368 12768 12374
rect 12714 12336 12716 12345
rect 12768 12336 12770 12345
rect 12714 12271 12770 12280
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11354 12204 11630
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12912 11286 12940 12378
rect 13004 12322 13032 12786
rect 13096 12782 13124 12922
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 13096 12442 13124 12718
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13004 12306 13124 12322
rect 13004 12300 13136 12306
rect 13004 12294 13084 12300
rect 13084 12242 13136 12248
rect 12992 11688 13044 11694
rect 12992 11630 13044 11636
rect 13004 11354 13032 11630
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11716 7274 11744 10406
rect 11900 9586 11928 10474
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11992 7954 12020 11154
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12636 10606 12664 11086
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12636 10266 12664 10542
rect 12728 10390 12940 10418
rect 12728 10266 12756 10390
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9110 12112 9318
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12176 8922 12204 9522
rect 12360 8974 12388 9522
rect 12544 9518 12572 10134
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12452 9364 12480 9454
rect 12636 9364 12664 10202
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12728 9586 12756 10066
rect 12820 9654 12848 10202
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12912 9382 12940 10390
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13004 9450 13032 9930
rect 13096 9518 13124 9998
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 12452 9336 12664 9364
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12084 8906 12204 8922
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12084 8900 12216 8906
rect 12084 8894 12164 8900
rect 12084 8090 12112 8894
rect 12164 8842 12216 8848
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12544 8022 12572 8570
rect 12636 8566 12664 8978
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12728 8362 12756 8978
rect 12912 8634 12940 9318
rect 13004 8974 13032 9386
rect 13096 9042 13124 9454
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8634 13124 8842
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 12544 7274 12572 7958
rect 13188 7954 13216 17070
rect 13372 16658 13400 17682
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13464 15162 13492 16050
rect 13556 15706 13584 17138
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13464 14550 13492 15098
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13648 11898 13676 17478
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13924 16658 13952 16934
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13728 16040 13780 16046
rect 13832 16028 13860 16390
rect 14016 16046 14044 17478
rect 14200 17134 14228 18566
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 17512 18222 17540 18566
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 15384 18148 15436 18154
rect 15384 18090 15436 18096
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 15396 17882 15424 18090
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 15384 17876 15436 17882
rect 15384 17818 15436 17824
rect 16684 17338 16712 18022
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 13780 16000 13860 16028
rect 14004 16040 14056 16046
rect 13728 15982 13780 15988
rect 14004 15982 14056 15988
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 14924 15700 14976 15706
rect 14924 15642 14976 15648
rect 14936 15026 14964 15642
rect 19076 15337 19104 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 19062 15328 19118 15337
rect 16900 15260 17208 15269
rect 19062 15263 19118 15272
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 14936 13938 14964 14962
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 13912 12708 13964 12714
rect 13832 12668 13912 12696
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13832 11014 13860 12668
rect 13912 12650 13964 12656
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14004 11620 14056 11626
rect 14004 11562 14056 11568
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10470 13860 10950
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13832 10062 13860 10406
rect 13924 10130 13952 11494
rect 14016 10674 14044 11562
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 15120 10470 15148 11698
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9178 13308 9862
rect 13832 9602 13860 9998
rect 15672 9926 15700 10542
rect 18604 10464 18656 10470
rect 18604 10406 18656 10412
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 13740 9574 13860 9602
rect 13740 9518 13768 9574
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13372 9042 13400 9454
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13372 8294 13400 8978
rect 13740 8974 13768 9454
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13832 9178 13860 9386
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 14108 9110 14136 9862
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12636 7342 12664 7686
rect 12728 7342 12756 7686
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12544 7002 12572 7210
rect 12820 7206 12848 7890
rect 13372 7886 13400 8230
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12912 7342 12940 7686
rect 13740 7410 13768 8910
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 13728 7404 13780 7410
rect 13728 7346 13780 7352
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 13188 6934 13216 7142
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13740 6866 13768 7346
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 8680 2746 8800 2774
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 8680 400 8708 2746
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 11164 400 11192 6122
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 13648 400 13676 5510
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 16132 400 16160 9862
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 18616 400 18644 10406
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
rect 11150 0 11206 400
rect 13634 0 13690 400
rect 16118 0 16174 400
rect 18602 0 18658 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 8758 13776 8814 13832
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 9218 10240 9274 10296
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 11058 12300 11114 12336
rect 11058 12280 11060 12300
rect 11060 12280 11112 12300
rect 11112 12280 11114 12300
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 12714 12316 12716 12336
rect 12716 12316 12768 12336
rect 12768 12316 12770 12336
rect 12714 12280 12770 12316
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 19062 15272 19118 15328
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 17902 15268 17908 15332
rect 17972 15330 17978 15332
rect 19057 15330 19123 15333
rect 17972 15328 19123 15330
rect 17972 15272 19062 15328
rect 19118 15272 19123 15328
rect 17972 15270 19123 15272
rect 17972 15268 17978 15270
rect 19057 15267 19123 15270
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 8753 13834 8819 13837
rect 8886 13834 8892 13836
rect 8753 13832 8892 13834
rect 8753 13776 8758 13832
rect 8814 13776 8892 13832
rect 8753 13774 8892 13776
rect 8753 13771 8819 13774
rect 8886 13772 8892 13774
rect 8956 13772 8962 13836
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 8886 12276 8892 12340
rect 8956 12338 8962 12340
rect 11053 12338 11119 12341
rect 8956 12336 11119 12338
rect 8956 12280 11058 12336
rect 11114 12280 11119 12336
rect 8956 12278 11119 12280
rect 8956 12276 8962 12278
rect 11053 12275 11119 12278
rect 12709 12338 12775 12341
rect 17902 12338 17908 12340
rect 12709 12336 17908 12338
rect 12709 12280 12714 12336
rect 12770 12280 17908 12336
rect 12709 12278 17908 12280
rect 12709 12275 12775 12278
rect 17902 12276 17908 12278
rect 17972 12276 17978 12340
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 8886 10236 8892 10300
rect 8956 10298 8962 10300
rect 9213 10298 9279 10301
rect 8956 10296 9279 10298
rect 8956 10240 9218 10296
rect 9274 10240 9279 10296
rect 8956 10238 9279 10240
rect 8956 10236 8962 10238
rect 9213 10235 9279 10238
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 16896 9759 17212 9760
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19253 8127 19569 8128
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 17908 15268 17972 15332
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 8892 13772 8956 13836
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 8892 12276 8956 12340
rect 17908 12276 17972 12340
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 8892 10236 8956 10300
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 8891 13836 8957 13837
rect 8891 13772 8892 13836
rect 8956 13772 8957 13836
rect 8891 13771 8957 13772
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 8894 12341 8954 13771
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 8891 12340 8957 12341
rect 8891 12276 8892 12340
rect 8956 12276 8957 12340
rect 8891 12275 8957 12276
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 8894 10301 8954 12275
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 8891 10300 8957 10301
rect 8891 10236 8892 10300
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 17907 15332 17973 15333
rect 17907 15268 17908 15332
rect 17972 15268 17973 15332
rect 17907 15267 17973 15268
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 17910 12341 17970 15267
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 17907 12340 17973 12341
rect 17907 12276 17908 12340
rect 17972 12276 17973 12340
rect 17907 12275 17973 12276
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__o221a_1  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9384 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10580 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8464 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11040 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9660 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9200 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _162_
timestamp 1704896540
transform 1 0 10212 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10488 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11316 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1704896540
transform -1 0 10488 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1704896540
transform 1 0 12604 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13984 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11040 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11316 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _172_
timestamp 1704896540
transform 1 0 11868 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _174_
timestamp 1704896540
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _175_
timestamp 1704896540
transform 1 0 11960 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _176_
timestamp 1704896540
transform -1 0 12788 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _177_
timestamp 1704896540
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12880 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _179_
timestamp 1704896540
transform -1 0 12788 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _180_
timestamp 1704896540
transform 1 0 12144 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1704896540
transform 1 0 11684 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1704896540
transform -1 0 13800 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13524 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13064 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _185_
timestamp 1704896540
transform -1 0 12880 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 1704896540
transform 1 0 13064 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1704896540
transform -1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1704896540
transform 1 0 6532 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _189_
timestamp 1704896540
transform -1 0 7360 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _190_
timestamp 1704896540
transform 1 0 6624 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _191_
timestamp 1704896540
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1704896540
transform 1 0 6072 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _193_
timestamp 1704896540
transform 1 0 5888 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _194_
timestamp 1704896540
transform -1 0 5704 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1704896540
transform 1 0 4968 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 1704896540
transform -1 0 7728 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _197_
timestamp 1704896540
transform 1 0 6532 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 1704896540
transform 1 0 6440 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _200_
timestamp 1704896540
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _201_
timestamp 1704896540
transform 1 0 4968 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1704896540
transform 1 0 11776 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _203_
timestamp 1704896540
transform 1 0 12788 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _204_
timestamp 1704896540
transform 1 0 12236 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1704896540
transform 1 0 12236 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _206_
timestamp 1704896540
transform -1 0 13248 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _207_
timestamp 1704896540
transform -1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _208_
timestamp 1704896540
transform 1 0 12144 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1704896540
transform -1 0 13064 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 1704896540
transform 1 0 12328 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp 1704896540
transform 1 0 12788 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _212_
timestamp 1704896540
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _213_
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _214_
timestamp 1704896540
transform -1 0 12144 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _215_
timestamp 1704896540
transform -1 0 10120 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _216_
timestamp 1704896540
transform -1 0 10396 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _217_
timestamp 1704896540
transform -1 0 10856 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1704896540
transform -1 0 10764 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _219_
timestamp 1704896540
transform 1 0 8556 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _220_
timestamp 1704896540
transform 1 0 9108 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _221_
timestamp 1704896540
transform -1 0 9660 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _222_
timestamp 1704896540
transform 1 0 6624 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _223_
timestamp 1704896540
transform 1 0 6072 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1704896540
transform -1 0 9292 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _225_
timestamp 1704896540
transform 1 0 5980 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _226_
timestamp 1704896540
transform -1 0 5704 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1704896540
transform 1 0 5060 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _228_
timestamp 1704896540
transform -1 0 6440 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _229_
timestamp 1704896540
transform 1 0 6716 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _230_
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1704896540
transform -1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp 1704896540
transform -1 0 8004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _233_
timestamp 1704896540
transform 1 0 7360 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _234_
timestamp 1704896540
transform 1 0 6900 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1704896540
transform -1 0 17204 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1704896540
transform 1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _238_
timestamp 1704896540
transform 1 0 12144 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13432 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _240_
timestamp 1704896540
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1704896540
transform -1 0 13984 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _242_
timestamp 1704896540
transform -1 0 13340 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _243_
timestamp 1704896540
transform 1 0 12696 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1704896540
transform 1 0 12420 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1704896540
transform 1 0 10856 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _246_
timestamp 1704896540
transform 1 0 11684 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1704896540
transform 1 0 11592 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _248_
timestamp 1704896540
transform 1 0 10120 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _249_
timestamp 1704896540
transform -1 0 11684 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1704896540
transform 1 0 9844 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _251_
timestamp 1704896540
transform -1 0 9292 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _252_
timestamp 1704896540
transform -1 0 9384 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1704896540
transform 1 0 9200 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _254_
timestamp 1704896540
transform 1 0 7820 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _255_
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1704896540
transform 1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _257_
timestamp 1704896540
transform -1 0 7452 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _258_
timestamp 1704896540
transform -1 0 6992 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1704896540
transform 1 0 7268 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _260_
timestamp 1704896540
transform -1 0 7176 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _261_
timestamp 1704896540
transform -1 0 6716 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7268 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _265_
timestamp 1704896540
transform 1 0 8556 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8648 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _267_
timestamp 1704896540
transform -1 0 11408 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _269_
timestamp 1704896540
transform -1 0 13248 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _270_
timestamp 1704896540
transform 1 0 9476 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _271_
timestamp 1704896540
transform 1 0 9568 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _272_
timestamp 1704896540
transform -1 0 10856 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _273_
timestamp 1704896540
transform 1 0 6440 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9476 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _277_
timestamp 1704896540
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1704896540
transform -1 0 13708 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _279_
timestamp 1704896540
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1704896540
transform -1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _282_
timestamp 1704896540
transform -1 0 8280 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 1704896540
transform 1 0 7544 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1704896540
transform 1 0 7084 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _285_
timestamp 1704896540
transform 1 0 9844 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1704896540
transform 1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1704896540
transform -1 0 7176 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1704896540
transform -1 0 13156 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _290_
timestamp 1704896540
transform 1 0 7268 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _291_
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1704896540
transform -1 0 11592 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _293_
timestamp 1704896540
transform 1 0 8188 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1704896540
transform 1 0 9936 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _296_
timestamp 1704896540
transform 1 0 8648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _297_
timestamp 1704896540
transform -1 0 8464 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _298_
timestamp 1704896540
transform 1 0 9384 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _299_
timestamp 1704896540
transform -1 0 10396 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _300_
timestamp 1704896540
transform -1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _301_
timestamp 1704896540
transform -1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _302_
timestamp 1704896540
transform 1 0 11500 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14996 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _304_
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _305_
timestamp 1704896540
transform 1 0 11040 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _306_
timestamp 1704896540
transform 1 0 9384 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _307_
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp 1704896540
transform 1 0 7360 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp 1704896540
transform 1 0 4784 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp 1704896540
transform 1 0 5428 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _312_
timestamp 1704896540
transform -1 0 6624 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _313_
timestamp 1704896540
transform -1 0 8188 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _314_
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _315_
timestamp 1704896540
transform 1 0 9292 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _316_
timestamp 1704896540
transform 1 0 9108 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _317_
timestamp 1704896540
transform 1 0 14076 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _318_
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _319_
timestamp 1704896540
transform -1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _320_
timestamp 1704896540
transform -1 0 13800 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _321_
timestamp 1704896540
transform 1 0 13708 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _322_
timestamp 1704896540
transform 1 0 13800 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _323_
timestamp 1704896540
transform -1 0 8096 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _324_
timestamp 1704896540
transform 1 0 4416 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _325_
timestamp 1704896540
transform 1 0 4048 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1704896540
transform 1 0 4140 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1704896540
transform -1 0 14996 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1704896540
transform -1 0 14996 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1704896540
transform -1 0 10488 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1704896540
transform 1 0 4232 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1704896540
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1704896540
transform -1 0 8280 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15088 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _335__12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15456 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12788 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 9292 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 8832 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 13248 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 12880 0 -1 15776
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1704896540
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_201
timestamp 1704896540
transform 1 0 19044 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18308 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp 1704896540
transform 1 0 19044 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1704896540
transform 1 0 19044 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 1704896540
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1704896540
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1704896540
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1704896540
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_201
timestamp 1704896540
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1704896540
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1704896540
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1704896540
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1704896540
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_201
timestamp 1704896540
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14260 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1704896540
transform 1 0 15364 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 15916 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_193
timestamp 1704896540
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_201
timestamp 1704896540
transform 1 0 19044 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_114
timestamp 1704896540
transform 1 0 11040 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_126
timestamp 1704896540
transform 1 0 12144 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1704896540
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1704896540
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1704896540
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1704896540
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1704896540
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1704896540
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1704896540
transform 1 0 6348 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_92
timestamp 1704896540
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12052 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_144
timestamp 1704896540
transform 1 0 13800 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1704896540
transform 1 0 14904 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17204 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_193
timestamp 1704896540
transform 1 0 18308 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_201
timestamp 1704896540
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_72
timestamp 1704896540
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1704896540
transform 1 0 8004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_104
timestamp 1704896540
transform 1 0 10120 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_112
timestamp 1704896540
transform 1 0 10856 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1704896540
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1704896540
transform 1 0 17940 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1704896540
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1704896540
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_86
timestamp 1704896540
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_101
timestamp 1704896540
transform 1 0 9844 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_122
timestamp 1704896540
transform 1 0 11776 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_133
timestamp 1704896540
transform 1 0 12788 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14260 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1704896540
transform 1 0 15364 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 15916 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_193
timestamp 1704896540
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_201
timestamp 1704896540
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_69
timestamp 1704896540
transform 1 0 6900 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1704896540
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_97
timestamp 1704896540
transform 1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_105
timestamp 1704896540
transform 1 0 10212 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_117
timestamp 1704896540
transform 1 0 11316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_125
timestamp 1704896540
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1704896540
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1704896540
transform 1 0 17940 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1704896540
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1704896540
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1704896540
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4140 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_47
timestamp 1704896540
transform 1 0 4876 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_75
timestamp 1704896540
transform 1 0 7452 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_87
timestamp 1704896540
transform 1 0 8556 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9108 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1704896540
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12052 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_160
timestamp 1704896540
transform 1 0 15272 0 -1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17204 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_193
timestamp 1704896540
transform 1 0 18308 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_201
timestamp 1704896540
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1704896540
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_114
timestamp 1704896540
transform 1 0 11040 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_120
timestamp 1704896540
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_159
timestamp 1704896540
transform 1 0 15180 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_171
timestamp 1704896540
transform 1 0 16284 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_183
timestamp 1704896540
transform 1 0 17388 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1704896540
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1704896540
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1704896540
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_70
timestamp 1704896540
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1704896540
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_116
timestamp 1704896540
transform 1 0 11224 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_128
timestamp 1704896540
transform 1 0 12328 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_144
timestamp 1704896540
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1704896540
transform 1 0 15824 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17204 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_193
timestamp 1704896540
transform 1 0 18308 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_201
timestamp 1704896540
transform 1 0 19044 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_65
timestamp 1704896540
transform 1 0 6532 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_69
timestamp 1704896540
transform 1 0 6900 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_74
timestamp 1704896540
transform 1 0 7360 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_78
timestamp 1704896540
transform 1 0 7728 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1704896540
transform 1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_105
timestamp 1704896540
transform 1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_117
timestamp 1704896540
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_123
timestamp 1704896540
transform 1 0 11868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1704896540
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_160
timestamp 1704896540
transform 1 0 15272 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_172
timestamp 1704896540
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_184
timestamp 1704896540
transform 1 0 17480 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1704896540
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1704896540
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5244 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_65
timestamp 1704896540
transform 1 0 6532 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_73
timestamp 1704896540
transform 1 0 7268 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9108 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_101
timestamp 1704896540
transform 1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_127
timestamp 1704896540
transform 1 0 12236 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_136
timestamp 1704896540
transform 1 0 13064 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_158
timestamp 1704896540
transform 1 0 15088 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1704896540
transform 1 0 15824 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1704896540
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_193
timestamp 1704896540
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp 1704896540
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1704896540
transform 1 0 3956 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_54
timestamp 1704896540
transform 1 0 5520 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_78
timestamp 1704896540
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_94
timestamp 1704896540
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_108
timestamp 1704896540
transform 1 0 10488 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_122
timestamp 1704896540
transform 1 0 11776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_132
timestamp 1704896540
transform 1 0 12696 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_146
timestamp 1704896540
transform 1 0 13984 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_158
timestamp 1704896540
transform 1 0 15088 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_170
timestamp 1704896540
transform 1 0 16192 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_182
timestamp 1704896540
transform 1 0 17296 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1704896540
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1704896540
transform 1 0 19044 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3036 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_73
timestamp 1704896540
transform 1 0 7268 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_80
timestamp 1704896540
transform 1 0 7912 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_92
timestamp 1704896540
transform 1 0 9016 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1704896540
transform 1 0 9384 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1704896540
transform 1 0 10580 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1704896540
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1704896540
transform 1 0 14260 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1704896540
transform 1 0 15364 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1704896540
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp 1704896540
transform 1 0 18308 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1704896540
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4324 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_47
timestamp 1704896540
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_69
timestamp 1704896540
transform 1 0 6900 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1704896540
transform 1 0 8004 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_105
timestamp 1704896540
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_121
timestamp 1704896540
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_136
timestamp 1704896540
transform 1 0 13064 0 1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_157
timestamp 1704896540
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_169
timestamp 1704896540
transform 1 0 16100 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_181
timestamp 1704896540
transform 1 0 17204 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1704896540
transform 1 0 18308 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1704896540
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4140 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5244 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_64
timestamp 1704896540
transform 1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_68
timestamp 1704896540
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_81
timestamp 1704896540
transform 1 0 8004 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_108
timestamp 1704896540
transform 1 0 10488 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_125
timestamp 1704896540
transform 1 0 12052 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1704896540
transform 1 0 13156 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1704896540
transform 1 0 14260 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15364 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 15916 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17204 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_193
timestamp 1704896540
transform 1 0 18308 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_201
timestamp 1704896540
transform 1 0 19044 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_57
timestamp 1704896540
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_88
timestamp 1704896540
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_104
timestamp 1704896540
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_116
timestamp 1704896540
transform 1 0 11224 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_120
timestamp 1704896540
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1704896540
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_157
timestamp 1704896540
transform 1 0 14996 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_169
timestamp 1704896540
transform 1 0 16100 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_181
timestamp 1704896540
transform 1 0 17204 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 1704896540
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_201
timestamp 1704896540
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4140 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_67
timestamp 1704896540
transform 1 0 6716 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_95
timestamp 1704896540
transform 1 0 9292 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_126
timestamp 1704896540
transform 1 0 12144 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_138
timestamp 1704896540
transform 1 0 13248 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_150
timestamp 1704896540
transform 1 0 14352 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_162
timestamp 1704896540
transform 1 0 15456 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_193
timestamp 1704896540
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_201
timestamp 1704896540
transform 1 0 19044 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 1932 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4324 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_52
timestamp 1704896540
transform 1 0 5336 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_66
timestamp 1704896540
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_78
timestamp 1704896540
transform 1 0 7728 0 1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_97
timestamp 1704896540
transform 1 0 9476 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_105
timestamp 1704896540
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_111
timestamp 1704896540
transform 1 0 10764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_123
timestamp 1704896540
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_131
timestamp 1704896540
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1704896540
transform 1 0 13064 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_157
timestamp 1704896540
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_169
timestamp 1704896540
transform 1 0 16100 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_181
timestamp 1704896540
transform 1 0 17204 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1704896540
transform 1 0 18308 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp 1704896540
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 828 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1704896540
transform 1 0 1932 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3036 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_39
timestamp 1704896540
transform 1 0 4140 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_57
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_63
timestamp 1704896540
transform 1 0 6348 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_72
timestamp 1704896540
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_80
timestamp 1704896540
transform 1 0 7912 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_86
timestamp 1704896540
transform 1 0 8464 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_94
timestamp 1704896540
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_129
timestamp 1704896540
transform 1 0 12420 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_133
timestamp 1704896540
transform 1 0 12788 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1704896540
transform 1 0 14720 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1704896540
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_193
timestamp 1704896540
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_201
timestamp 1704896540
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 1932 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_53
timestamp 1704896540
transform 1 0 5428 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1704896540
transform 1 0 8004 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_106
timestamp 1704896540
transform 1 0 10304 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_110
timestamp 1704896540
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_118
timestamp 1704896540
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_126
timestamp 1704896540
transform 1 0 12144 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1704896540
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_148
timestamp 1704896540
transform 1 0 14168 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_160
timestamp 1704896540
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_172
timestamp 1704896540
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_184
timestamp 1704896540
transform 1 0 17480 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1704896540
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1704896540
transform 1 0 1932 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1704896540
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1704896540
transform 1 0 5244 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1704896540
transform 1 0 5796 0 -1 16864
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_73
timestamp 1704896540
transform 1 0 7268 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_85
timestamp 1704896540
transform 1 0 8372 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_97
timestamp 1704896540
transform 1 0 9476 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_109
timestamp 1704896540
transform 1 0 10580 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_125
timestamp 1704896540
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_133
timestamp 1704896540
transform 1 0 12788 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_139
timestamp 1704896540
transform 1 0 13340 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_146
timestamp 1704896540
transform 1 0 13984 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_158
timestamp 1704896540
transform 1 0 15088 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1704896540
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp 1704896540
transform 1 0 18308 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1704896540
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3036 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4324 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_45
timestamp 1704896540
transform 1 0 4692 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_75
timestamp 1704896540
transform 1 0 7452 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_96
timestamp 1704896540
transform 1 0 9384 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_109
timestamp 1704896540
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_123
timestamp 1704896540
transform 1 0 11868 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_130
timestamp 1704896540
transform 1 0 12512 0 1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_157
timestamp 1704896540
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_169
timestamp 1704896540
transform 1 0 16100 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_181
timestamp 1704896540
transform 1 0 17204 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_193
timestamp 1704896540
transform 1 0 18308 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1704896540
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1704896540
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1704896540
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1704896540
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1704896540
transform 1 0 5244 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1704896540
transform 1 0 5612 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_57
timestamp 1704896540
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_72
timestamp 1704896540
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_95
timestamp 1704896540
transform 1 0 9292 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_132
timestamp 1704896540
transform 1 0 12696 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_146
timestamp 1704896540
transform 1 0 13984 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_158
timestamp 1704896540
transform 1 0 15088 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1704896540
transform 1 0 15732 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1704896540
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1704896540
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp 1704896540
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_201
timestamp 1704896540
transform 1 0 19044 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1704896540
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_76
timestamp 1704896540
transform 1 0 7544 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_104
timestamp 1704896540
transform 1 0 10120 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_112
timestamp 1704896540
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_130
timestamp 1704896540
transform 1 0 12512 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_157
timestamp 1704896540
transform 1 0 14996 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_181
timestamp 1704896540
transform 1 0 17204 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_193
timestamp 1704896540
transform 1 0 18308 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1704896540
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_14
timestamp 1704896540
transform 1 0 1840 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_25
timestamp 1704896540
transform 1 0 2852 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_29
timestamp 1704896540
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_37
timestamp 1704896540
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp 1704896540
transform 1 0 4508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1704896540
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_61
timestamp 1704896540
transform 1 0 6164 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_73
timestamp 1704896540
transform 1 0 7268 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_79
timestamp 1704896540
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp 1704896540
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_85
timestamp 1704896540
transform 1 0 8372 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_99
timestamp 1704896540
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1704896540
transform 1 0 10764 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_116
timestamp 1704896540
transform 1 0 11224 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_128
timestamp 1704896540
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_133
timestamp 1704896540
transform 1 0 12788 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1704896540
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_141
timestamp 1704896540
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_147
timestamp 1704896540
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1704896540
transform 1 0 14444 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1704896540
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1704896540
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_172
timestamp 1704896540
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_187
timestamp 1704896540
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1704896540
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1704896540
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1704896540
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6440 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 6532 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 5888 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 7268 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 7268 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 11040 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16376 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 14444 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform -1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1704896540
transform 1 0 2576 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 920 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1704896540
transform 1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1704896540
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1704896540
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1704896540
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1704896540
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 10061 19040 10061 19040 4 VGND
rlabel metal1 s 9982 18496 9982 18496 4 VPWR
rlabel metal1 s 16843 18122 16843 18122 4 _000_
rlabel metal1 s 14034 18122 14034 18122 4 _001_
rlabel metal1 s 13600 17034 13600 17034 4 _002_
rlabel metal2 s 12374 17986 12374 17986 4 _003_
rlabel metal1 s 10345 17714 10345 17714 4 _004_
rlabel metal2 s 8689 18190 8689 18190 4 _005_
rlabel metal2 s 9062 17510 9062 17510 4 _006_
rlabel metal1 s 5699 17034 5699 17034 4 _007_
rlabel metal2 s 6026 17986 6026 17986 4 _008_
rlabel metal1 s 7544 11186 7544 11186 4 _009_
rlabel metal2 s 6302 7548 6302 7548 4 _010_
rlabel metal2 s 7866 7276 7866 7276 4 _011_
rlabel metal2 s 8694 7548 8694 7548 4 _012_
rlabel metal2 s 9614 7922 9614 7922 4 _013_
rlabel metal1 s 9338 6834 9338 6834 4 _014_
rlabel metal1 s 14168 10098 14168 10098 4 _015_
rlabel metal1 s 13938 10642 13938 10642 4 _016_
rlabel metal1 s 11642 7310 11642 7310 4 _017_
rlabel metal1 s 13344 6902 13344 6902 4 _018_
rlabel metal1 s 13800 9146 13800 9146 4 _019_
rlabel metal2 s 14117 9078 14117 9078 4 _020_
rlabel metal1 s 7452 9146 7452 9146 4 _021_
rlabel metal1 s 4968 9146 4968 9146 4 _022_
rlabel metal1 s 5796 11322 5796 11322 4 _023_
rlabel metal1 s 4733 12342 4733 12342 4 _024_
rlabel metal1 s 13416 12682 13416 12682 4 _025_
rlabel metal1 s 13850 14858 13850 14858 4 _026_
rlabel metal1 s 13942 13838 13942 13838 4 _027_
rlabel metal1 s 10902 15130 10902 15130 4 _028_
rlabel metal1 s 9940 13430 9940 13430 4 _029_
rlabel metal2 s 5106 15334 5106 15334 4 _030_
rlabel metal1 s 5331 13838 5331 13838 4 _031_
rlabel metal2 s 7682 13634 7682 13634 4 _032_
rlabel metal1 s 7268 17510 7268 17510 4 _033_
rlabel metal1 s 6716 17850 6716 17850 4 _034_
rlabel metal2 s 7406 15742 7406 15742 4 _035_
rlabel metal1 s 7452 15402 7452 15402 4 _036_
rlabel metal2 s 9062 15810 9062 15810 4 _037_
rlabel metal2 s 9154 15810 9154 15810 4 _038_
rlabel metal2 s 9246 16218 9246 16218 4 _039_
rlabel metal2 s 10534 15708 10534 15708 4 _040_
rlabel metal1 s 13386 16014 13386 16014 4 _041_
rlabel metal2 s 12466 15742 12466 15742 4 _042_
rlabel metal1 s 10120 15402 10120 15402 4 _043_
rlabel metal1 s 10166 15504 10166 15504 4 _044_
rlabel metal1 s 10074 15334 10074 15334 4 _045_
rlabel metal1 s 6716 15674 6716 15674 4 _046_
rlabel metal1 s 8786 16048 8786 16048 4 _047_
rlabel metal1 s 10120 12750 10120 12750 4 _048_
rlabel metal1 s 9614 14348 9614 14348 4 _049_
rlabel metal1 s 12742 13362 12742 13362 4 _050_
rlabel metal1 s 13616 17510 13616 17510 4 _051_
rlabel metal2 s 6670 14756 6670 14756 4 _052_
rlabel metal2 s 8142 12070 8142 12070 4 _053_
rlabel metal2 s 12650 9962 12650 9962 4 _054_
rlabel metal2 s 8050 12036 8050 12036 4 _055_
rlabel metal1 s 9706 12614 9706 12614 4 _056_
rlabel metal1 s 8878 12750 8878 12750 4 _057_
rlabel metal2 s 6302 8092 6302 8092 4 _058_
rlabel metal1 s 12926 7990 12926 7990 4 _059_
rlabel metal1 s 7866 7514 7866 7514 4 _060_
rlabel metal1 s 12190 7752 12190 7752 4 _061_
rlabel metal1 s 6026 7854 6026 7854 4 _062_
rlabel metal1 s 11408 16966 11408 16966 4 _063_
rlabel metal2 s 8970 7514 8970 7514 4 _064_
rlabel metal1 s 11040 7854 11040 7854 4 _065_
rlabel metal1 s 8418 8024 8418 8024 4 _066_
rlabel metal1 s 8602 6698 8602 6698 4 _067_
rlabel metal1 s 10304 9010 10304 9010 4 _068_
rlabel metal1 s 10350 9146 10350 9146 4 _069_
rlabel metal2 s 9154 8092 9154 8092 4 _070_
rlabel metal2 s 9062 9996 9062 9996 4 _071_
rlabel metal1 s 12466 7276 12466 7276 4 _072_
rlabel metal1 s 9062 9588 9062 9588 4 _073_
rlabel metal1 s 9660 9010 9660 9010 4 _074_
rlabel metal1 s 9798 9418 9798 9418 4 _075_
rlabel metal1 s 10488 9622 10488 9622 4 _076_
rlabel metal1 s 9384 16966 9384 16966 4 _077_
rlabel metal2 s 8970 9724 8970 9724 4 _078_
rlabel metal2 s 9430 9180 9430 9180 4 _079_
rlabel metal2 s 10718 10132 10718 10132 4 _080_
rlabel metal1 s 11040 11118 11040 11118 4 _081_
rlabel metal2 s 11086 10982 11086 10982 4 _082_
rlabel metal2 s 10810 11458 10810 11458 4 _083_
rlabel metal1 s 12627 11186 12627 11186 4 _084_
rlabel metal2 s 13018 11492 13018 11492 4 _085_
rlabel metal1 s 12098 11696 12098 11696 4 _086_
rlabel metal1 s 12190 11152 12190 11152 4 _087_
rlabel metal1 s 12144 11322 12144 11322 4 _088_
rlabel metal1 s 11040 8058 11040 8058 4 _089_
rlabel metal2 s 12650 7514 12650 7514 4 _090_
rlabel metal2 s 12742 7514 12742 7514 4 _091_
rlabel metal1 s 12926 9656 12926 9656 4 _092_
rlabel metal2 s 12650 8772 12650 8772 4 _093_
rlabel metal1 s 12052 9146 12052 9146 4 _094_
rlabel metal1 s 13570 9044 13570 9044 4 _095_
rlabel metal1 s 13386 9146 13386 9146 4 _096_
rlabel metal2 s 12558 9826 12558 9826 4 _097_
rlabel metal2 s 12834 9928 12834 9928 4 _098_
rlabel metal1 s 13524 10098 13524 10098 4 _099_
rlabel metal1 s 6854 9044 6854 9044 4 _100_
rlabel metal1 s 6946 8976 6946 8976 4 _101_
rlabel metal2 s 5842 9248 5842 9248 4 _102_
rlabel metal2 s 6678 12614 6678 12614 4 _103_
rlabel metal1 s 5750 9146 5750 9146 4 _104_
rlabel metal1 s 5106 9010 5106 9010 4 _105_
rlabel metal1 s 5980 12614 5980 12614 4 _106_
rlabel metal2 s 6302 11356 6302 11356 4 _107_
rlabel metal1 s 12650 12852 12650 12852 4 _108_
rlabel metal1 s 5520 12750 5520 12750 4 _109_
rlabel metal1 s 12466 12784 12466 12784 4 _110_
rlabel metal1 s 12696 12138 12696 12138 4 _111_
rlabel metal2 s 12282 14858 12282 14858 4 _112_
rlabel metal1 s 12834 14348 12834 14348 4 _113_
rlabel metal1 s 12236 14042 12236 14042 4 _114_
rlabel metal1 s 12696 14926 12696 14926 4 _115_
rlabel metal1 s 12696 13498 12696 13498 4 _116_
rlabel metal1 s 12788 13226 12788 13226 4 _117_
rlabel metal1 s 10810 14246 10810 14246 4 _118_
rlabel metal1 s 9890 13872 9890 13872 4 _119_
rlabel metal1 s 9154 14484 9154 14484 4 _120_
rlabel metal1 s 10350 14552 10350 14552 4 _121_
rlabel metal2 s 10442 14756 10442 14756 4 _122_
rlabel metal1 s 9430 12784 9430 12784 4 _123_
rlabel metal2 s 9154 13396 9154 13396 4 _124_
rlabel metal1 s 7176 14790 7176 14790 4 _125_
rlabel metal1 s 5796 14246 5796 14246 4 _126_
rlabel metal1 s 6302 14382 6302 14382 4 _127_
rlabel metal1 s 5796 14314 5796 14314 4 _128_
rlabel metal1 s 5290 14348 5290 14348 4 _129_
rlabel metal1 s 6302 13498 6302 13498 4 _130_
rlabel metal2 s 7314 14042 7314 14042 4 _131_
rlabel metal2 s 7130 13702 7130 13702 4 _132_
rlabel metal2 s 7866 14246 7866 14246 4 _133_
rlabel metal1 s 7314 13362 7314 13362 4 _134_
rlabel metal1 s 13202 17714 13202 17714 4 _135_
rlabel metal1 s 13938 17510 13938 17510 4 _136_
rlabel metal2 s 13386 17170 13386 17170 4 _137_
rlabel metal1 s 12880 17850 12880 17850 4 _138_
rlabel metal1 s 13570 16422 13570 16422 4 _139_
rlabel metal2 s 12926 16864 12926 16864 4 _140_
rlabel metal1 s 12604 17510 12604 17510 4 _141_
rlabel metal1 s 11500 17306 11500 17306 4 _142_
rlabel metal2 s 10350 17170 10350 17170 4 _143_
rlabel metal2 s 10534 17442 10534 17442 4 _144_
rlabel metal2 s 9246 17782 9246 17782 4 _145_
rlabel metal1 s 9108 17850 9108 17850 4 _146_
rlabel metal1 s 9154 16762 9154 16762 4 _147_
rlabel metal1 s 8326 16966 8326 16966 4 _148_
rlabel metal1 s 7452 16626 7452 16626 4 _149_
rlabel metal1 s 6992 16966 6992 16966 4 _150_
rlabel metal3 s 18515 15300 18515 15300 4 clk
rlabel metal1 s 13110 11254 13110 11254 4 clknet_0_clk
rlabel metal1 s 4324 9554 4324 9554 4 clknet_2_0__leaf_clk
rlabel metal1 s 4278 13838 4278 13838 4 clknet_2_1__leaf_clk
rlabel metal1 s 13754 12750 13754 12750 4 clknet_2_2__leaf_clk
rlabel metal1 s 13294 17170 13294 17170 4 clknet_2_3__leaf_clk
rlabel metal1 s 13386 9520 13386 9520 4 counter\[0\]
rlabel metal2 s 12466 14552 12466 14552 4 counter\[10\]
rlabel metal1 s 11086 16082 11086 16082 4 counter\[11\]
rlabel metal2 s 8602 15708 8602 15708 4 counter\[12\]
rlabel metal2 s 8878 16014 8878 16014 4 counter\[13\]
rlabel metal1 s 6836 16014 6836 16014 4 counter\[14\]
rlabel metal2 s 7038 16252 7038 16252 4 counter\[15\]
rlabel metal2 s 12558 7480 12558 7480 4 counter\[1\]
rlabel metal1 s 12834 10064 12834 10064 4 counter\[2\]
rlabel metal1 s 13018 8874 13018 8874 4 counter\[3\]
rlabel metal1 s 6118 9486 6118 9486 4 counter\[4\]
rlabel metal1 s 5980 9690 5980 9690 4 counter\[5\]
rlabel metal1 s 6762 12954 6762 12954 4 counter\[6\]
rlabel metal1 s 6394 12716 6394 12716 4 counter\[7\]
rlabel metal2 s 13018 15062 13018 15062 4 counter\[8\]
rlabel metal1 s 13386 16082 13386 16082 4 counter\[9\]
rlabel metal1 s 16054 18802 16054 18802 4 data[0]
rlabel metal1 s 14260 18802 14260 18802 4 data[1]
rlabel metal1 s 12604 18802 12604 18802 4 data[2]
rlabel metal1 s 10902 18802 10902 18802 4 data[3]
rlabel metal1 s 9384 18802 9384 18802 4 data[4]
rlabel metal1 s 7544 18802 7544 18802 4 data[5]
rlabel metal1 s 5888 18802 5888 18802 4 data[6]
rlabel metal1 s 4232 18802 4232 18802 4 data[7]
rlabel metal2 s 13754 17884 13754 17884 4 divider\[0\]
rlabel metal2 s 13938 16796 13938 16796 4 divider\[1\]
rlabel metal2 s 12466 17884 12466 17884 4 divider\[2\]
rlabel metal2 s 11638 17306 11638 17306 4 divider\[3\]
rlabel metal1 s 9844 18190 9844 18190 4 divider\[4\]
rlabel metal2 s 8694 17068 8694 17068 4 divider\[5\]
rlabel metal2 s 6394 16796 6394 16796 4 divider\[6\]
rlabel metal1 s 7314 18224 7314 18224 4 divider\[7\]
rlabel metal1 s 2576 18802 2576 18802 4 ext_data
rlabel metal1 s 920 18802 920 18802 4 load_divider
rlabel metal1 s 17572 18802 17572 18802 4 n_rst
rlabel metal2 s 13202 18428 13202 18428 4 net1
rlabel metal2 s 6946 18462 6946 18462 4 net10
rlabel metal1 s 17342 18190 17342 18190 4 net11
rlabel metal1 s 15456 17850 15456 17850 4 net12
rlabel metal1 s 5290 12784 5290 12784 4 net13
rlabel metal2 s 6118 11356 6118 11356 4 net14
rlabel metal2 s 7222 9214 7222 9214 4 net15
rlabel metal1 s 6532 7922 6532 7922 4 net16
rlabel metal2 s 8694 7004 8694 7004 4 net17
rlabel metal1 s 10120 8602 10120 8602 4 net18
rlabel metal1 s 13708 17102 13708 17102 4 net2
rlabel metal2 s 12558 18122 12558 18122 4 net3
rlabel metal1 s 11040 17646 11040 17646 4 net4
rlabel metal1 s 8878 18700 8878 18700 4 net5
rlabel metal1 s 8740 17170 8740 17170 4 net6
rlabel metal1 s 6578 17170 6578 17170 4 net7
rlabel metal1 s 6118 17714 6118 17714 4 net8
rlabel metal2 s 6302 17340 6302 17340 4 net9
rlabel metal2 s 1242 1860 1242 1860 4 r2r_out[0]
rlabel metal1 s 4324 7242 4324 7242 4 r2r_out[1]
rlabel metal1 s 6394 6630 6394 6630 4 r2r_out[2]
rlabel metal2 s 8694 1557 8694 1557 4 r2r_out[3]
rlabel metal1 s 11086 6154 11086 6154 4 r2r_out[4]
rlabel metal2 s 13662 2948 13662 2948 4 r2r_out[5]
rlabel metal1 s 15916 9894 15916 9894 4 r2r_out[6]
rlabel metal1 s 16882 10438 16882 10438 4 r2r_out[7]
rlabel metal2 s 16698 17680 16698 17680 4 rst
flabel metal4 s 19251 496 19571 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14536 496 14856 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9821 496 10141 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5106 496 5426 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16894 496 17214 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12179 496 12499 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7464 496 7784 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2749 496 3069 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 19062 19600 19118 20000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 15750 19600 15806 20000 0 FreeSans 280 90 0 0 data[0]
port 4 nsew
flabel metal2 s 14094 19600 14150 20000 0 FreeSans 280 90 0 0 data[1]
port 5 nsew
flabel metal2 s 12438 19600 12494 20000 0 FreeSans 280 90 0 0 data[2]
port 6 nsew
flabel metal2 s 10782 19600 10838 20000 0 FreeSans 280 90 0 0 data[3]
port 7 nsew
flabel metal2 s 9126 19600 9182 20000 0 FreeSans 280 90 0 0 data[4]
port 8 nsew
flabel metal2 s 7470 19600 7526 20000 0 FreeSans 280 90 0 0 data[5]
port 9 nsew
flabel metal2 s 5814 19600 5870 20000 0 FreeSans 280 90 0 0 data[6]
port 10 nsew
flabel metal2 s 4158 19600 4214 20000 0 FreeSans 280 90 0 0 data[7]
port 11 nsew
flabel metal2 s 2502 19600 2558 20000 0 FreeSans 280 90 0 0 ext_data
port 12 nsew
flabel metal2 s 846 19600 902 20000 0 FreeSans 280 90 0 0 load_divider
port 13 nsew
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 280 90 0 0 n_rst
port 14 nsew
flabel metal2 s 1214 0 1270 400 0 FreeSans 280 90 0 0 r2r_out[0]
port 15 nsew
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 r2r_out[1]
port 16 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 r2r_out[2]
port 17 nsew
flabel metal2 s 8666 0 8722 400 0 FreeSans 280 90 0 0 r2r_out[3]
port 18 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 r2r_out[4]
port 19 nsew
flabel metal2 s 13634 0 13690 400 0 FreeSans 280 90 0 0 r2r_out[5]
port 20 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 r2r_out[6]
port 21 nsew
flabel metal2 s 18602 0 18658 400 0 FreeSans 280 90 0 0 r2r_out[7]
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string GDS_END 930526
string GDS_FILE ../gds/r2r_dac_control.gds
string GDS_START 281042
<< end >>
