** sch_path: /home/matt/work/asic-workshop/shuttle-tt08/tt08-analog-r2r-dac-3v3/xschem/r2r.sch
.subckt r2r b4 b2 b1 b0 b5 b6 b7 b3 out VGND
*.PININFO b0:I b1:I b2:I b3:I b4:I b5:I b6:I b7:I out:O VGND:B
XR1 net1 b0 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR7 net2 b1 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR10 net3 b2 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR13 net4 b3 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR16 net5 b4 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR19 net6 b5 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR22 net7 b6 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR25 net8 b7 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR5 b a VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR8 c b VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR11 d c VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR14 e d VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR17 f e VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR20 g f VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR23 out g VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR3 net9 a VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR2 a net1 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR6 b net2 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR9 c net3 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR12 d net4 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR15 e net5 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR18 f net6 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR21 g net7 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR24 out net8 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR4 VGND net9 VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR26 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
XR27 VGND VGND VGND sky130_fd_pr__res_high_po_1p41 L=45 mult=1 m=1
.ends
.end
