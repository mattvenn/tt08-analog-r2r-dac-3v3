magic
tech sky130A
magscale 1 2
timestamp 1720442423
<< viali >>
rect 2789 18921 2823 18955
rect 949 18785 983 18819
rect 2605 18785 2639 18819
rect 4261 18785 4295 18819
rect 5917 18785 5951 18819
rect 7573 18785 7607 18819
rect 9229 18785 9263 18819
rect 11161 18785 11195 18819
rect 12725 18785 12759 18819
rect 14381 18785 14415 18819
rect 16313 18785 16347 18819
rect 17693 18785 17727 18819
rect 1225 18717 1259 18751
rect 4445 18649 4479 18683
rect 6101 18581 6135 18615
rect 7757 18581 7791 18615
rect 9413 18581 9447 18615
rect 10977 18581 11011 18615
rect 12541 18581 12575 18615
rect 14197 18581 14231 18615
rect 16129 18581 16163 18615
rect 17509 18581 17543 18615
rect 7481 18377 7515 18411
rect 10057 18309 10091 18343
rect 7205 18241 7239 18275
rect 4353 18173 4387 18207
rect 7573 18173 7607 18207
rect 7665 18173 7699 18207
rect 8401 18173 8435 18207
rect 9873 18173 9907 18207
rect 10241 18173 10275 18207
rect 10425 18173 10459 18207
rect 17049 18173 17083 18207
rect 4620 18105 4654 18139
rect 6960 18105 6994 18139
rect 8668 18105 8702 18139
rect 5733 18037 5767 18071
rect 5825 18037 5859 18071
rect 7297 18037 7331 18071
rect 9781 18037 9815 18071
rect 10241 18037 10275 18071
rect 15853 18037 15887 18071
rect 16957 18037 16991 18071
rect 6929 17833 6963 17867
rect 7021 17833 7055 17867
rect 7665 17833 7699 17867
rect 8125 17833 8159 17867
rect 8217 17833 8251 17867
rect 8861 17833 8895 17867
rect 16405 17765 16439 17799
rect 4077 17697 4111 17731
rect 4344 17697 4378 17731
rect 6561 17697 6595 17731
rect 6745 17697 6779 17731
rect 7389 17697 7423 17731
rect 7757 17697 7791 17731
rect 8585 17697 8619 17731
rect 8677 17697 8711 17731
rect 8953 17697 8987 17731
rect 9680 17697 9714 17731
rect 10977 17697 11011 17731
rect 6469 17629 6503 17663
rect 7481 17629 7515 17663
rect 7849 17629 7883 17663
rect 9045 17629 9079 17663
rect 9413 17629 9447 17663
rect 16129 17629 16163 17663
rect 5457 17561 5491 17595
rect 10793 17561 10827 17595
rect 5825 17493 5859 17527
rect 6745 17493 6779 17527
rect 7941 17493 7975 17527
rect 9137 17493 9171 17527
rect 9321 17493 9355 17527
rect 11069 17493 11103 17527
rect 17877 17493 17911 17527
rect 4077 17289 4111 17323
rect 6929 17289 6963 17323
rect 8769 17289 8803 17323
rect 11345 17289 11379 17323
rect 6101 17221 6135 17255
rect 4445 17153 4479 17187
rect 7113 17153 7147 17187
rect 7573 17153 7607 17187
rect 9505 17153 9539 17187
rect 9873 17153 9907 17187
rect 9965 17153 9999 17187
rect 2329 17085 2363 17119
rect 2513 17085 2547 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4629 17085 4663 17119
rect 4721 17085 4755 17119
rect 6009 17085 6043 17119
rect 6285 17085 6319 17119
rect 7205 17085 7239 17119
rect 8861 17085 8895 17119
rect 10149 17085 10183 17119
rect 10241 17085 10275 17119
rect 10425 17085 10459 17119
rect 4445 17017 4479 17051
rect 11253 17017 11287 17051
rect 2421 16949 2455 16983
rect 6377 16949 6411 16983
rect 10333 16949 10367 16983
rect 9505 16745 9539 16779
rect 2320 16677 2354 16711
rect 3709 16677 3743 16711
rect 3985 16609 4019 16643
rect 4169 16609 4203 16643
rect 4436 16609 4470 16643
rect 9689 16609 9723 16643
rect 10057 16609 10091 16643
rect 2053 16541 2087 16575
rect 3709 16541 3743 16575
rect 6377 16541 6411 16575
rect 3433 16473 3467 16507
rect 5549 16473 5583 16507
rect 3893 16405 3927 16439
rect 5825 16405 5859 16439
rect 9965 16405 9999 16439
rect 3709 16201 3743 16235
rect 4721 16201 4755 16235
rect 10517 16201 10551 16235
rect 13185 16201 13219 16235
rect 4537 16133 4571 16167
rect 4997 16133 5031 16167
rect 12633 16133 12667 16167
rect 2053 16065 2087 16099
rect 5825 16065 5859 16099
rect 6101 16065 6135 16099
rect 7113 16065 7147 16099
rect 13553 16065 13587 16099
rect 1409 15997 1443 16031
rect 1777 15997 1811 16031
rect 1869 15997 1903 16031
rect 3433 15997 3467 16031
rect 3617 15997 3651 16031
rect 4353 15997 4387 16031
rect 5181 15997 5215 16031
rect 5365 15997 5399 16031
rect 5733 15997 5767 16031
rect 7225 15997 7259 16031
rect 7389 15997 7423 16031
rect 7573 15997 7607 16031
rect 7665 15997 7699 16031
rect 7757 15997 7791 16031
rect 7941 15997 7975 16031
rect 9137 15997 9171 16031
rect 11069 15997 11103 16031
rect 11345 15997 11379 16031
rect 13829 15997 13863 16031
rect 14381 15997 14415 16031
rect 14565 15997 14599 16031
rect 4705 15929 4739 15963
rect 4905 15929 4939 15963
rect 6837 15929 6871 15963
rect 7021 15929 7055 15963
rect 7113 15929 7147 15963
rect 9382 15929 9416 15963
rect 13001 15929 13035 15963
rect 13921 15929 13955 15963
rect 14197 15929 14231 15963
rect 1685 15861 1719 15895
rect 2605 15861 2639 15895
rect 3249 15861 3283 15895
rect 8125 15861 8159 15895
rect 13201 15861 13235 15895
rect 13369 15861 13403 15895
rect 13737 15861 13771 15895
rect 14105 15861 14139 15895
rect 3709 15657 3743 15691
rect 4629 15657 4663 15691
rect 7205 15657 7239 15691
rect 7573 15657 7607 15691
rect 9229 15657 9263 15691
rect 9873 15657 9907 15691
rect 11345 15657 11379 15691
rect 12817 15657 12851 15691
rect 4169 15589 4203 15623
rect 1970 15521 2004 15555
rect 2237 15521 2271 15555
rect 3249 15521 3283 15555
rect 3341 15521 3375 15555
rect 3525 15521 3559 15555
rect 4445 15521 4479 15555
rect 4537 15521 4571 15555
rect 4721 15521 4755 15555
rect 6653 15521 6687 15555
rect 6929 15521 6963 15555
rect 7021 15521 7055 15555
rect 7456 15521 7490 15555
rect 8033 15521 8067 15555
rect 8217 15521 8251 15555
rect 8309 15521 8343 15555
rect 8401 15521 8435 15555
rect 8677 15521 8711 15555
rect 9413 15521 9447 15555
rect 9505 15521 9539 15555
rect 11529 15521 11563 15555
rect 11805 15521 11839 15555
rect 11989 15521 12023 15555
rect 12449 15521 12483 15555
rect 12541 15521 12575 15555
rect 12725 15521 12759 15555
rect 12909 15521 12943 15555
rect 13645 15521 13679 15555
rect 13912 15521 13946 15555
rect 15209 15521 15243 15555
rect 2789 15453 2823 15487
rect 2881 15453 2915 15487
rect 2973 15453 3007 15487
rect 3065 15453 3099 15487
rect 4169 15453 4203 15487
rect 7665 15453 7699 15487
rect 7941 15453 7975 15487
rect 8769 15453 8803 15487
rect 12265 15453 12299 15487
rect 12357 15453 12391 15487
rect 13093 15453 13127 15487
rect 13185 15453 13219 15487
rect 13277 15453 13311 15487
rect 13369 15453 13403 15487
rect 6745 15385 6779 15419
rect 8585 15385 8619 15419
rect 857 15317 891 15351
rect 2605 15317 2639 15351
rect 4353 15317 4387 15351
rect 7297 15317 7331 15351
rect 8677 15317 8711 15351
rect 9045 15317 9079 15351
rect 12081 15317 12115 15351
rect 13553 15317 13587 15351
rect 15025 15317 15059 15351
rect 15393 15317 15427 15351
rect 2421 15113 2455 15147
rect 2881 15113 2915 15147
rect 11161 15113 11195 15147
rect 11529 15113 11563 15147
rect 12817 15113 12851 15147
rect 16865 15113 16899 15147
rect 2053 15045 2087 15079
rect 2697 15045 2731 15079
rect 14151 15045 14185 15079
rect 4905 14977 4939 15011
rect 11897 14977 11931 15011
rect 13093 14977 13127 15011
rect 13277 14977 13311 15011
rect 15117 14977 15151 15011
rect 15393 14977 15427 15011
rect 6653 14909 6687 14943
rect 9965 14909 9999 14943
rect 10701 14909 10735 14943
rect 10977 14909 11011 14943
rect 11161 14909 11195 14943
rect 11713 14909 11747 14943
rect 13001 14909 13035 14943
rect 13185 14909 13219 14943
rect 13553 14909 13587 14943
rect 13737 14909 13771 14943
rect 13921 14909 13955 14943
rect 16865 14909 16899 14943
rect 16957 14909 16991 14943
rect 2421 14841 2455 14875
rect 3065 14841 3099 14875
rect 5089 14841 5123 14875
rect 8217 14841 8251 14875
rect 9698 14841 9732 14875
rect 10793 14841 10827 14875
rect 2605 14773 2639 14807
rect 2865 14773 2899 14807
rect 8585 14773 8619 14807
rect 13553 14773 13587 14807
rect 16681 14773 16715 14807
rect 17233 14773 17267 14807
rect 6837 14569 6871 14603
rect 7757 14569 7791 14603
rect 8033 14569 8067 14603
rect 8861 14569 8895 14603
rect 9505 14569 9539 14603
rect 13461 14569 13495 14603
rect 16773 14569 16807 14603
rect 4721 14501 4755 14535
rect 6193 14501 6227 14535
rect 1961 14433 1995 14467
rect 2228 14433 2262 14467
rect 3985 14433 4019 14467
rect 4169 14433 4203 14467
rect 4261 14433 4295 14467
rect 4445 14433 4479 14467
rect 5181 14433 5215 14467
rect 5365 14433 5399 14467
rect 6469 14433 6503 14467
rect 6745 14433 6779 14467
rect 7021 14433 7055 14467
rect 7205 14433 7239 14467
rect 7573 14433 7607 14467
rect 8125 14433 8159 14467
rect 9321 14433 9355 14467
rect 11529 14433 11563 14467
rect 13369 14433 13403 14467
rect 13553 14433 13587 14467
rect 15025 14433 15059 14467
rect 15301 14433 15335 14467
rect 16497 14433 16531 14467
rect 16957 14433 16991 14467
rect 17141 14433 17175 14467
rect 17233 14433 17267 14467
rect 4353 14365 4387 14399
rect 5089 14365 5123 14399
rect 7297 14365 7331 14399
rect 7389 14365 7423 14399
rect 9229 14365 9263 14399
rect 11253 14365 11287 14399
rect 12173 14365 12207 14399
rect 4077 14297 4111 14331
rect 5825 14297 5859 14331
rect 6377 14297 6411 14331
rect 11437 14297 11471 14331
rect 3341 14229 3375 14263
rect 4537 14229 4571 14263
rect 4721 14229 4755 14263
rect 5549 14229 5583 14263
rect 6193 14229 6227 14263
rect 6653 14229 6687 14263
rect 11345 14229 11379 14263
rect 11621 14229 11655 14263
rect 15117 14229 15151 14263
rect 15485 14229 15519 14263
rect 17233 14229 17267 14263
rect 17417 14229 17451 14263
rect 2053 14025 2087 14059
rect 5457 14025 5491 14059
rect 7757 14025 7791 14059
rect 13553 14025 13587 14059
rect 15117 14025 15151 14059
rect 16589 14025 16623 14059
rect 2421 13957 2455 13991
rect 5365 13957 5399 13991
rect 2329 13889 2363 13923
rect 6377 13889 6411 13923
rect 16773 13889 16807 13923
rect 17509 13889 17543 13923
rect 2237 13821 2271 13855
rect 2513 13821 2547 13855
rect 2605 13821 2639 13855
rect 2697 13821 2731 13855
rect 2881 13821 2915 13855
rect 3985 13821 4019 13855
rect 5641 13821 5675 13855
rect 5733 13821 5767 13855
rect 6644 13821 6678 13855
rect 11161 13821 11195 13855
rect 11417 13821 11451 13855
rect 12725 13821 12759 13855
rect 13369 13821 13403 13855
rect 13553 13821 13587 13855
rect 13829 13821 13863 13855
rect 14841 13821 14875 13855
rect 14933 13821 14967 13855
rect 15209 13821 15243 13855
rect 15476 13821 15510 13855
rect 4252 13753 4286 13787
rect 6009 13753 6043 13787
rect 15117 13753 15151 13787
rect 2789 13685 2823 13719
rect 5825 13685 5859 13719
rect 12541 13685 12575 13719
rect 13737 13685 13771 13719
rect 1501 13481 1535 13515
rect 2881 13481 2915 13515
rect 4445 13481 4479 13515
rect 18153 13481 18187 13515
rect 1133 13413 1167 13447
rect 1961 13413 1995 13447
rect 10333 13413 10367 13447
rect 11222 13413 11256 13447
rect 12541 13413 12575 13447
rect 12741 13413 12775 13447
rect 15761 13413 15795 13447
rect 857 13345 891 13379
rect 1041 13345 1075 13379
rect 1409 13345 1443 13379
rect 1685 13345 1719 13379
rect 4629 13345 4663 13379
rect 6745 13345 6779 13379
rect 6929 13345 6963 13379
rect 8493 13345 8527 13379
rect 8585 13345 8619 13379
rect 9045 13345 9079 13379
rect 9781 13345 9815 13379
rect 10517 13345 10551 13379
rect 10793 13345 10827 13379
rect 13921 13345 13955 13379
rect 14177 13345 14211 13379
rect 15485 13345 15519 13379
rect 16957 13345 16991 13379
rect 17509 13345 17543 13379
rect 18521 13345 18555 13379
rect 1133 13277 1167 13311
rect 1317 13277 1351 13311
rect 1869 13277 1903 13311
rect 2513 13277 2547 13311
rect 3433 13277 3467 13311
rect 8125 13277 8159 13311
rect 9137 13277 9171 13311
rect 9505 13277 9539 13311
rect 10977 13277 11011 13311
rect 13001 13277 13035 13311
rect 13277 13277 13311 13311
rect 18613 13277 18647 13311
rect 12909 13209 12943 13243
rect 15301 13209 15335 13243
rect 1041 13141 1075 13175
rect 6837 13141 6871 13175
rect 8769 13141 8803 13175
rect 8861 13141 8895 13175
rect 9965 13141 9999 13175
rect 10701 13141 10735 13175
rect 12357 13141 12391 13175
rect 12725 13141 12759 13175
rect 16129 13141 16163 13175
rect 18797 13141 18831 13175
rect 3249 12937 3283 12971
rect 8033 12937 8067 12971
rect 8217 12937 8251 12971
rect 10977 12937 11011 12971
rect 13093 12937 13127 12971
rect 14013 12937 14047 12971
rect 18429 12937 18463 12971
rect 3709 12869 3743 12903
rect 13277 12869 13311 12903
rect 1041 12801 1075 12835
rect 3341 12801 3375 12835
rect 7941 12801 7975 12835
rect 12909 12801 12943 12835
rect 14473 12801 14507 12835
rect 14749 12801 14783 12835
rect 17049 12801 17083 12835
rect 3065 12733 3099 12767
rect 3525 12733 3559 12767
rect 7113 12733 7147 12767
rect 7665 12733 7699 12767
rect 8493 12733 8527 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 11621 12733 11655 12767
rect 11805 12733 11839 12767
rect 12081 12733 12115 12767
rect 12265 12733 12299 12767
rect 12357 12733 12391 12767
rect 12725 12733 12759 12767
rect 13093 12733 13127 12767
rect 13553 12733 13587 12767
rect 13829 12733 13863 12767
rect 13921 12733 13955 12767
rect 14381 12733 14415 12767
rect 16129 12733 16163 12767
rect 17316 12733 17350 12767
rect 2820 12665 2854 12699
rect 3249 12665 3283 12699
rect 8760 12665 8794 12699
rect 12817 12665 12851 12699
rect 13645 12665 13679 12699
rect 16773 12665 16807 12699
rect 1593 12597 1627 12631
rect 1685 12597 1719 12631
rect 5825 12597 5859 12631
rect 9873 12597 9907 12631
rect 11161 12597 11195 12631
rect 11621 12597 11655 12631
rect 12449 12597 12483 12631
rect 12633 12597 12667 12631
rect 857 12393 891 12427
rect 4077 12393 4111 12427
rect 4921 12393 4955 12427
rect 6837 12393 6871 12427
rect 9597 12393 9631 12427
rect 1970 12325 2004 12359
rect 2421 12325 2455 12359
rect 2621 12325 2655 12359
rect 4721 12325 4755 12359
rect 6929 12325 6963 12359
rect 7389 12325 7423 12359
rect 12357 12325 12391 12359
rect 13921 12325 13955 12359
rect 3985 12257 4019 12291
rect 4169 12257 4203 12291
rect 4261 12257 4295 12291
rect 5365 12257 5399 12291
rect 5549 12257 5583 12291
rect 6469 12257 6503 12291
rect 7021 12257 7055 12291
rect 7205 12257 7239 12291
rect 7297 12257 7331 12291
rect 8686 12257 8720 12291
rect 8953 12257 8987 12291
rect 9045 12257 9079 12291
rect 9321 12257 9355 12291
rect 11069 12257 11103 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 17325 12257 17359 12291
rect 17509 12257 17543 12291
rect 2237 12189 2271 12223
rect 6561 12189 6595 12223
rect 11253 12189 11287 12223
rect 11621 12189 11655 12223
rect 12173 12189 12207 12223
rect 5181 12121 5215 12155
rect 2605 12053 2639 12087
rect 2789 12053 2823 12087
rect 4445 12053 4479 12087
rect 4905 12053 4939 12087
rect 5089 12053 5123 12087
rect 7573 12053 7607 12087
rect 9229 12053 9263 12087
rect 11437 12053 11471 12087
rect 16497 12053 16531 12087
rect 2881 11849 2915 11883
rect 4537 11849 4571 11883
rect 5089 11849 5123 11883
rect 7021 11849 7055 11883
rect 9505 11849 9539 11883
rect 12357 11849 12391 11883
rect 14289 11849 14323 11883
rect 15209 11849 15243 11883
rect 3985 11781 4019 11815
rect 4629 11781 4663 11815
rect 2697 11713 2731 11747
rect 3249 11713 3283 11747
rect 4997 11713 5031 11747
rect 6469 11713 6503 11747
rect 13185 11713 13219 11747
rect 14473 11713 14507 11747
rect 2973 11645 3007 11679
rect 3893 11645 3927 11679
rect 4169 11645 4203 11679
rect 4261 11645 4295 11679
rect 6653 11645 6687 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 11152 11645 11186 11679
rect 12541 11645 12575 11679
rect 12725 11645 12759 11679
rect 12909 11645 12943 11679
rect 13093 11645 13127 11679
rect 13553 11645 13587 11679
rect 14013 11645 14047 11679
rect 14381 11645 14415 11679
rect 14565 11645 14599 11679
rect 15025 11645 15059 11679
rect 15117 11645 15151 11679
rect 16313 11645 16347 11679
rect 16773 11645 16807 11679
rect 2697 11577 2731 11611
rect 3985 11577 4019 11611
rect 6202 11577 6236 11611
rect 6837 11577 6871 11611
rect 13737 11577 13771 11611
rect 14105 11577 14139 11611
rect 14289 11577 14323 11611
rect 12265 11509 12299 11543
rect 13921 11509 13955 11543
rect 15393 11509 15427 11543
rect 15945 11509 15979 11543
rect 3433 11305 3467 11339
rect 5641 11305 5675 11339
rect 6009 11305 6043 11339
rect 2053 11169 2087 11203
rect 2320 11169 2354 11203
rect 4261 11169 4295 11203
rect 4528 11169 4562 11203
rect 5825 11169 5859 11203
rect 8769 11169 8803 11203
rect 8953 11169 8987 11203
rect 9137 11169 9171 11203
rect 9321 11169 9355 11203
rect 9413 11169 9447 11203
rect 9597 11169 9631 11203
rect 12633 11169 12667 11203
rect 13277 11169 13311 11203
rect 14841 11169 14875 11203
rect 16589 11169 16623 11203
rect 17141 11169 17175 11203
rect 17693 11169 17727 11203
rect 14105 11101 14139 11135
rect 14933 11101 14967 11135
rect 16681 11101 16715 11135
rect 8861 11033 8895 11067
rect 9229 11033 9263 11067
rect 9505 11033 9539 11067
rect 16957 10965 16991 10999
rect 10793 10693 10827 10727
rect 10149 10625 10183 10659
rect 12633 10625 12667 10659
rect 8401 10557 8435 10591
rect 8585 10557 8619 10591
rect 10057 10557 10091 10591
rect 10609 10557 10643 10591
rect 10793 10557 10827 10591
rect 12725 10557 12759 10591
rect 14105 10557 14139 10591
rect 14289 10557 14323 10591
rect 14565 10557 14599 10591
rect 14841 10557 14875 10591
rect 16405 10557 16439 10591
rect 16589 10557 16623 10591
rect 17049 10557 17083 10591
rect 14381 10489 14415 10523
rect 14933 10489 14967 10523
rect 18061 10489 18095 10523
rect 8493 10421 8527 10455
rect 13369 10421 13403 10455
rect 14197 10421 14231 10455
rect 14749 10421 14783 10455
rect 16681 10217 16715 10251
rect 9873 10149 9907 10183
rect 15209 10149 15243 10183
rect 16313 10149 16347 10183
rect 9689 10081 9723 10115
rect 10287 10081 10321 10115
rect 10425 10081 10459 10115
rect 10517 10081 10551 10115
rect 10609 10081 10643 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 11253 10081 11287 10115
rect 11345 10081 11379 10115
rect 13829 10081 13863 10115
rect 14013 10081 14047 10115
rect 14289 10081 14323 10115
rect 14565 10081 14599 10115
rect 14749 10081 14783 10115
rect 15025 10081 15059 10115
rect 15301 10081 15335 10115
rect 16497 10081 16531 10115
rect 16773 10081 16807 10115
rect 17417 10081 17451 10115
rect 10149 10013 10183 10047
rect 14473 10013 14507 10047
rect 14841 10013 14875 10047
rect 10057 9945 10091 9979
rect 14381 9945 14415 9979
rect 17233 9945 17267 9979
rect 10793 9877 10827 9911
rect 11621 9877 11655 9911
rect 13921 9877 13955 9911
rect 14105 9877 14139 9911
rect 13001 9673 13035 9707
rect 8861 9605 8895 9639
rect 10609 9605 10643 9639
rect 13553 9605 13587 9639
rect 16405 9605 16439 9639
rect 9689 9537 9723 9571
rect 10425 9537 10459 9571
rect 11897 9537 11931 9571
rect 12173 9537 12207 9571
rect 12817 9537 12851 9571
rect 13737 9537 13771 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 8861 9469 8895 9503
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 9597 9469 9631 9503
rect 10885 9469 10919 9503
rect 12081 9469 12115 9503
rect 12265 9469 12299 9503
rect 12357 9469 12391 9503
rect 13093 9469 13127 9503
rect 13185 9469 13219 9503
rect 13369 9469 13403 9503
rect 13829 9469 13863 9503
rect 14381 9469 14415 9503
rect 15853 9469 15887 9503
rect 16037 9469 16071 9503
rect 10241 9401 10275 9435
rect 10609 9401 10643 9435
rect 14565 9401 14599 9435
rect 15945 9401 15979 9435
rect 9229 9333 9263 9367
rect 9781 9333 9815 9367
rect 10149 9333 10183 9367
rect 10793 9333 10827 9367
rect 12541 9333 12575 9367
rect 13185 9333 13219 9367
rect 14197 9333 14231 9367
rect 16773 9333 16807 9367
rect 10149 9129 10183 9163
rect 12909 9129 12943 9163
rect 13645 9129 13679 9163
rect 15485 9129 15519 9163
rect 16589 9129 16623 9163
rect 17509 9129 17543 9163
rect 11069 9061 11103 9095
rect 9229 8993 9263 9027
rect 10057 8993 10091 9027
rect 13093 8993 13127 9027
rect 13185 8993 13219 9027
rect 13829 8993 13863 9027
rect 14565 8993 14599 9027
rect 14657 8993 14691 9027
rect 14749 8993 14783 9027
rect 14933 8993 14967 9027
rect 15669 8993 15703 9027
rect 15853 8993 15887 9027
rect 15945 8993 15979 9027
rect 16497 8993 16531 9027
rect 16957 8993 16991 9027
rect 17601 8993 17635 9027
rect 17693 8993 17727 9027
rect 17877 8993 17911 9027
rect 17969 8993 18003 9027
rect 18245 8993 18279 9027
rect 18429 8993 18463 9027
rect 9505 8925 9539 8959
rect 13277 8925 13311 8959
rect 13369 8925 13403 8959
rect 13921 8925 13955 8959
rect 14013 8925 14047 8959
rect 14105 8925 14139 8959
rect 16681 8925 16715 8959
rect 17233 8925 17267 8959
rect 12357 8857 12391 8891
rect 14289 8857 14323 8891
rect 18245 8857 18279 8891
rect 7941 8789 7975 8823
rect 16129 8789 16163 8823
rect 17049 8789 17083 8823
rect 18153 8789 18187 8823
rect 11805 8585 11839 8619
rect 12909 8585 12943 8619
rect 15393 8585 15427 8619
rect 16589 8585 16623 8619
rect 8493 8517 8527 8551
rect 12725 8517 12759 8551
rect 14657 8517 14691 8551
rect 16957 8517 16991 8551
rect 9873 8449 9907 8483
rect 11621 8449 11655 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 15853 8449 15887 8483
rect 16681 8449 16715 8483
rect 18153 8449 18187 8483
rect 9606 8381 9640 8415
rect 11897 8381 11931 8415
rect 12173 8381 12207 8415
rect 12265 8381 12299 8415
rect 13553 8381 13587 8415
rect 14013 8381 14047 8415
rect 14197 8381 14231 8415
rect 14289 8381 14323 8415
rect 14381 8381 14415 8415
rect 14933 8381 14967 8415
rect 15025 8381 15059 8415
rect 15209 8381 15243 8415
rect 15301 8381 15335 8415
rect 15393 8381 15427 8415
rect 15577 8381 15611 8415
rect 15669 8381 15703 8415
rect 15945 8381 15979 8415
rect 16589 8381 16623 8415
rect 17233 8381 17267 8415
rect 17509 8381 17543 8415
rect 17969 8381 18003 8415
rect 11621 8313 11655 8347
rect 12877 8313 12911 8347
rect 13093 8313 13127 8347
rect 13737 8313 13771 8347
rect 13921 8313 13955 8347
rect 14749 8313 14783 8347
rect 17049 8313 17083 8347
rect 11989 8245 12023 8279
rect 12449 8245 12483 8279
rect 17417 8245 17451 8279
rect 17601 8245 17635 8279
rect 18061 8245 18095 8279
rect 9965 8041 9999 8075
rect 11345 8041 11379 8075
rect 12173 8041 12207 8075
rect 13277 8041 13311 8075
rect 14657 8041 14691 8075
rect 17877 8041 17911 8075
rect 9781 7973 9815 8007
rect 11437 7973 11471 8007
rect 12909 7973 12943 8007
rect 15301 7973 15335 8007
rect 15531 7939 15565 7973
rect 10057 7905 10091 7939
rect 12449 7905 12483 7939
rect 12541 7905 12575 7939
rect 12633 7905 12667 7939
rect 12817 7905 12851 7939
rect 13093 7905 13127 7939
rect 13369 7905 13403 7939
rect 13737 7905 13771 7939
rect 14473 7905 14507 7939
rect 14657 7905 14691 7939
rect 17049 7905 17083 7939
rect 17233 7905 17267 7939
rect 17325 7905 17359 7939
rect 17417 7905 17451 7939
rect 17785 7905 17819 7939
rect 17969 7905 18003 7939
rect 18061 7905 18095 7939
rect 18245 7905 18279 7939
rect 11621 7837 11655 7871
rect 10977 7769 11011 7803
rect 9781 7701 9815 7735
rect 13553 7701 13587 7735
rect 15485 7701 15519 7735
rect 15669 7701 15703 7735
rect 17693 7701 17727 7735
rect 18061 7701 18095 7735
rect 17417 7497 17451 7531
rect 10057 7361 10091 7395
rect 11069 7361 11103 7395
rect 11253 7361 11287 7395
rect 12265 7361 12299 7395
rect 17509 7361 17543 7395
rect 9781 7293 9815 7327
rect 10977 7293 11011 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 13921 7293 13955 7327
rect 14105 7293 14139 7327
rect 14197 7293 14231 7327
rect 14289 7293 14323 7327
rect 14473 7293 14507 7327
rect 15025 7293 15059 7327
rect 16037 7293 16071 7327
rect 16313 7293 16347 7327
rect 17233 7293 17267 7327
rect 8401 7225 8435 7259
rect 12633 7225 12667 7259
rect 14381 7225 14415 7259
rect 15209 7225 15243 7259
rect 17049 7225 17083 7259
rect 10609 7157 10643 7191
rect 13737 7157 13771 7191
rect 15393 7157 15427 7191
rect 15853 7157 15887 7191
rect 16221 7157 16255 7191
rect 10057 6953 10091 6987
rect 11437 6953 11471 6987
rect 14657 6953 14691 6987
rect 16881 6953 16915 6987
rect 9965 6885 9999 6919
rect 11345 6885 11379 6919
rect 13277 6885 13311 6919
rect 16681 6885 16715 6919
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 9045 6817 9079 6851
rect 9137 6817 9171 6851
rect 9321 6817 9355 6851
rect 9413 6817 9447 6851
rect 10517 6817 10551 6851
rect 10609 6817 10643 6851
rect 10793 6817 10827 6851
rect 12173 6817 12207 6851
rect 12357 6817 12391 6851
rect 12909 6817 12943 6851
rect 13737 6817 13771 6851
rect 14013 6817 14047 6851
rect 14381 6817 14415 6851
rect 14654 6817 14688 6851
rect 15117 6817 15151 6851
rect 15485 6817 15519 6851
rect 15577 6817 15611 6851
rect 15669 6817 15703 6851
rect 10241 6749 10275 6783
rect 11621 6749 11655 6783
rect 11989 6749 12023 6783
rect 12265 6749 12299 6783
rect 12449 6749 12483 6783
rect 12817 6749 12851 6783
rect 13185 6749 13219 6783
rect 13829 6749 13863 6783
rect 15393 6749 15427 6783
rect 8769 6681 8803 6715
rect 9597 6681 9631 6715
rect 10793 6681 10827 6715
rect 12633 6681 12667 6715
rect 13921 6681 13955 6715
rect 14289 6681 14323 6715
rect 9137 6613 9171 6647
rect 10977 6613 11011 6647
rect 13553 6613 13587 6647
rect 14473 6613 14507 6647
rect 15025 6613 15059 6647
rect 15209 6613 15243 6647
rect 16865 6613 16899 6647
rect 17049 6613 17083 6647
rect 9689 6409 9723 6443
rect 14381 6409 14415 6443
rect 15117 6409 15151 6443
rect 16957 6409 16991 6443
rect 11069 6341 11103 6375
rect 14933 6341 14967 6375
rect 16773 6341 16807 6375
rect 17233 6341 17267 6375
rect 10149 6273 10183 6307
rect 10333 6273 10367 6307
rect 15301 6273 15335 6307
rect 15393 6273 15427 6307
rect 15577 6273 15611 6307
rect 16313 6273 16347 6307
rect 17141 6273 17175 6307
rect 10057 6205 10091 6239
rect 10793 6205 10827 6239
rect 11069 6205 11103 6239
rect 13829 6205 13863 6239
rect 14013 6205 14047 6239
rect 14197 6205 14231 6239
rect 14841 6205 14875 6239
rect 15025 6205 15059 6239
rect 15485 6205 15519 6239
rect 16405 6205 16439 6239
rect 16865 6205 16899 6239
rect 17233 6205 17267 6239
rect 17509 6205 17543 6239
rect 10885 6137 10919 6171
rect 14105 6137 14139 6171
rect 17141 6069 17175 6103
rect 17417 6069 17451 6103
rect 11590 5797 11624 5831
rect 9790 5729 9824 5763
rect 10057 5729 10091 5763
rect 11345 5729 11379 5763
rect 8677 5525 8711 5559
rect 12725 5525 12759 5559
rect 9413 5185 9447 5219
rect 10977 5185 11011 5219
rect 9680 5117 9714 5151
rect 16681 5117 16715 5151
rect 11244 5049 11278 5083
rect 16926 5049 16960 5083
rect 10793 4981 10827 5015
rect 12357 4981 12391 5015
rect 18061 4981 18095 5015
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 2777 18955 2835 18961
rect 2777 18921 2789 18955
rect 2823 18952 2835 18955
rect 10502 18952 10508 18964
rect 2823 18924 10508 18952
rect 2823 18921 2835 18924
rect 2777 18915 2835 18921
rect 10502 18912 10508 18924
rect 10560 18912 10566 18964
rect 842 18776 848 18828
rect 900 18816 906 18828
rect 937 18819 995 18825
rect 937 18816 949 18819
rect 900 18788 949 18816
rect 900 18776 906 18788
rect 937 18785 949 18788
rect 983 18785 995 18819
rect 937 18779 995 18785
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 2593 18819 2651 18825
rect 2593 18816 2605 18819
rect 2556 18788 2605 18816
rect 2556 18776 2562 18788
rect 2593 18785 2605 18788
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4212 18788 4261 18816
rect 4212 18776 4218 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5868 18788 5917 18816
rect 5868 18776 5874 18788
rect 5905 18785 5917 18788
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7524 18788 7573 18816
rect 7524 18776 7530 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 7561 18779 7619 18785
rect 9122 18776 9128 18828
rect 9180 18816 9186 18828
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 9180 18788 9229 18816
rect 9180 18776 9186 18788
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 11112 18788 11161 18816
rect 11112 18776 11118 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12492 18788 12725 18816
rect 12492 18776 12498 18788
rect 12713 18785 12725 18788
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14148 18788 14381 18816
rect 14148 18776 14154 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15804 18788 16313 18816
rect 15804 18776 15810 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17460 18788 17693 18816
rect 17460 18776 17466 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 1213 18751 1271 18757
rect 1213 18717 1225 18751
rect 1259 18748 1271 18751
rect 7190 18748 7196 18760
rect 1259 18720 7196 18748
rect 1259 18717 1271 18720
rect 1213 18711 1271 18717
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 4433 18683 4491 18689
rect 4433 18649 4445 18683
rect 4479 18680 4491 18683
rect 8018 18680 8024 18692
rect 4479 18652 8024 18680
rect 4479 18649 4491 18652
rect 4433 18643 4491 18649
rect 8018 18640 8024 18652
rect 8076 18640 8082 18692
rect 6089 18615 6147 18621
rect 6089 18581 6101 18615
rect 6135 18612 6147 18615
rect 6914 18612 6920 18624
rect 6135 18584 6920 18612
rect 6135 18581 6147 18584
rect 6089 18575 6147 18581
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 7745 18615 7803 18621
rect 7745 18581 7757 18615
rect 7791 18612 7803 18615
rect 8662 18612 8668 18624
rect 7791 18584 8668 18612
rect 7791 18581 7803 18584
rect 7745 18575 7803 18581
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 9398 18572 9404 18624
rect 9456 18572 9462 18624
rect 10226 18572 10232 18624
rect 10284 18612 10290 18624
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10284 18584 10977 18612
rect 10284 18572 10290 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 12618 18612 12624 18624
rect 12575 18584 12624 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 14182 18572 14188 18624
rect 14240 18572 14246 18624
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 16117 18615 16175 18621
rect 16117 18612 16129 18615
rect 15252 18584 16129 18612
rect 15252 18572 15258 18584
rect 16117 18581 16129 18584
rect 16163 18581 16175 18615
rect 16117 18575 16175 18581
rect 17494 18572 17500 18624
rect 17552 18572 17558 18624
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 7006 18368 7012 18420
rect 7064 18408 7070 18420
rect 7469 18411 7527 18417
rect 7469 18408 7481 18411
rect 7064 18380 7481 18408
rect 7064 18368 7070 18380
rect 7469 18377 7481 18380
rect 7515 18377 7527 18411
rect 7469 18371 7527 18377
rect 10045 18343 10103 18349
rect 10045 18309 10057 18343
rect 10091 18340 10103 18343
rect 10410 18340 10416 18352
rect 10091 18312 10416 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 10410 18300 10416 18312
rect 10468 18300 10474 18352
rect 7193 18275 7251 18281
rect 7193 18241 7205 18275
rect 7239 18272 7251 18275
rect 7239 18244 8432 18272
rect 7239 18241 7251 18244
rect 7193 18235 7251 18241
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4341 18207 4399 18213
rect 4341 18204 4353 18207
rect 4212 18176 4353 18204
rect 4212 18164 4218 18176
rect 4341 18173 4353 18176
rect 4387 18204 4399 18207
rect 7208 18204 7236 18235
rect 4387 18176 7236 18204
rect 4387 18173 4399 18176
rect 4341 18167 4399 18173
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7558 18204 7564 18216
rect 7340 18176 7564 18204
rect 7340 18164 7346 18176
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 8404 18213 8432 18244
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 9122 18204 9128 18216
rect 8435 18176 9128 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 4608 18139 4666 18145
rect 4608 18105 4620 18139
rect 4654 18136 4666 18139
rect 6948 18139 7006 18145
rect 4654 18108 6868 18136
rect 4654 18105 4666 18108
rect 4608 18099 4666 18105
rect 5718 18028 5724 18080
rect 5776 18028 5782 18080
rect 5813 18071 5871 18077
rect 5813 18037 5825 18071
rect 5859 18068 5871 18071
rect 6270 18068 6276 18080
rect 5859 18040 6276 18068
rect 5859 18037 5871 18040
rect 5813 18031 5871 18037
rect 6270 18028 6276 18040
rect 6328 18028 6334 18080
rect 6840 18068 6868 18108
rect 6948 18105 6960 18139
rect 6994 18136 7006 18139
rect 7466 18136 7472 18148
rect 6994 18108 7472 18136
rect 6994 18105 7006 18108
rect 6948 18099 7006 18105
rect 7466 18096 7472 18108
rect 7524 18096 7530 18148
rect 7098 18068 7104 18080
rect 6840 18040 7104 18068
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7282 18028 7288 18080
rect 7340 18028 7346 18080
rect 7374 18028 7380 18080
rect 7432 18068 7438 18080
rect 7668 18068 7696 18167
rect 9122 18164 9128 18176
rect 9180 18164 9186 18216
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9732 18176 9873 18204
rect 9732 18164 9738 18176
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 9861 18167 9919 18173
rect 10226 18164 10232 18216
rect 10284 18164 10290 18216
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10502 18204 10508 18216
rect 10459 18176 10508 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 10502 18164 10508 18176
rect 10560 18164 10566 18216
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 17494 18204 17500 18216
rect 17083 18176 17500 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 17494 18164 17500 18176
rect 17552 18164 17558 18216
rect 8656 18139 8714 18145
rect 8656 18105 8668 18139
rect 8702 18136 8714 18139
rect 8846 18136 8852 18148
rect 8702 18108 8852 18136
rect 8702 18105 8714 18108
rect 8656 18099 8714 18105
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 7742 18068 7748 18080
rect 7432 18040 7748 18068
rect 7432 18028 7438 18040
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 9674 18028 9680 18080
rect 9732 18068 9738 18080
rect 9769 18071 9827 18077
rect 9769 18068 9781 18071
rect 9732 18040 9781 18068
rect 9732 18028 9738 18040
rect 9769 18037 9781 18040
rect 9815 18037 9827 18071
rect 9769 18031 9827 18037
rect 10226 18028 10232 18080
rect 10284 18028 10290 18080
rect 15838 18028 15844 18080
rect 15896 18028 15902 18080
rect 16942 18028 16948 18080
rect 17000 18028 17006 18080
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 6917 17867 6975 17873
rect 6917 17833 6929 17867
rect 6963 17864 6975 17867
rect 7009 17867 7067 17873
rect 7009 17864 7021 17867
rect 6963 17836 7021 17864
rect 6963 17833 6975 17836
rect 6917 17827 6975 17833
rect 7009 17833 7021 17836
rect 7055 17833 7067 17867
rect 7374 17864 7380 17876
rect 7009 17827 7067 17833
rect 7208 17836 7380 17864
rect 7208 17796 7236 17836
rect 7374 17824 7380 17836
rect 7432 17824 7438 17876
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7524 17836 7665 17864
rect 7524 17824 7530 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 8113 17867 8171 17873
rect 8113 17833 8125 17867
rect 8159 17864 8171 17867
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 8159 17836 8217 17864
rect 8159 17833 8171 17836
rect 8113 17827 8171 17833
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 8205 17827 8263 17833
rect 8846 17824 8852 17876
rect 8904 17824 8910 17876
rect 10410 17796 10416 17808
rect 6564 17768 7236 17796
rect 7484 17768 10416 17796
rect 4065 17731 4123 17737
rect 4065 17697 4077 17731
rect 4111 17728 4123 17731
rect 4154 17728 4160 17740
rect 4111 17700 4160 17728
rect 4111 17697 4123 17700
rect 4065 17691 4123 17697
rect 4154 17688 4160 17700
rect 4212 17688 4218 17740
rect 4338 17737 4344 17740
rect 4332 17691 4344 17737
rect 4338 17688 4344 17691
rect 4396 17688 4402 17740
rect 6564 17737 6592 17768
rect 6549 17731 6607 17737
rect 6549 17697 6561 17731
rect 6595 17697 6607 17731
rect 6549 17691 6607 17697
rect 6733 17731 6791 17737
rect 6733 17697 6745 17731
rect 6779 17728 6791 17731
rect 7190 17728 7196 17740
rect 6779 17700 7196 17728
rect 6779 17697 6791 17700
rect 6733 17691 6791 17697
rect 7190 17688 7196 17700
rect 7248 17688 7254 17740
rect 7377 17734 7435 17737
rect 7484 17734 7512 17768
rect 8588 17740 8616 17768
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 15838 17756 15844 17808
rect 15896 17796 15902 17808
rect 16393 17799 16451 17805
rect 16393 17796 16405 17799
rect 15896 17768 16405 17796
rect 15896 17756 15902 17768
rect 16393 17765 16405 17768
rect 16439 17765 16451 17799
rect 16393 17759 16451 17765
rect 16942 17756 16948 17808
rect 17000 17756 17006 17808
rect 7377 17731 7512 17734
rect 7377 17697 7389 17731
rect 7423 17706 7512 17731
rect 7423 17697 7435 17706
rect 7377 17691 7435 17697
rect 7742 17688 7748 17740
rect 7800 17688 7806 17740
rect 8570 17688 8576 17740
rect 8628 17688 8634 17740
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 8938 17688 8944 17740
rect 8996 17688 9002 17740
rect 9490 17728 9496 17740
rect 9048 17700 9496 17728
rect 6454 17660 6460 17672
rect 5460 17632 6460 17660
rect 5460 17604 5488 17632
rect 6454 17620 6460 17632
rect 6512 17620 6518 17672
rect 7466 17620 7472 17672
rect 7524 17620 7530 17672
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 9048 17669 9076 17700
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 9668 17731 9726 17737
rect 9668 17697 9680 17731
rect 9714 17728 9726 17731
rect 10134 17728 10140 17740
rect 9714 17700 10140 17728
rect 9714 17697 9726 17700
rect 9668 17691 9726 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10796 17700 10977 17728
rect 7837 17663 7895 17669
rect 7837 17660 7849 17663
rect 7616 17632 7849 17660
rect 7616 17620 7622 17632
rect 7837 17629 7849 17632
rect 7883 17660 7895 17663
rect 9033 17663 9091 17669
rect 9033 17660 9045 17663
rect 7883 17632 9045 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 9033 17629 9045 17632
rect 9079 17629 9091 17663
rect 9033 17623 9091 17629
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9180 17632 9413 17660
rect 9180 17620 9186 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9401 17623 9459 17629
rect 5442 17552 5448 17604
rect 5500 17552 5506 17604
rect 6914 17552 6920 17604
rect 6972 17592 6978 17604
rect 6972 17564 7512 17592
rect 6972 17552 6978 17564
rect 7484 17536 7512 17564
rect 7742 17552 7748 17604
rect 7800 17592 7806 17604
rect 8938 17592 8944 17604
rect 7800 17564 8944 17592
rect 7800 17552 7806 17564
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 10796 17601 10824 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 15286 17620 15292 17672
rect 15344 17660 15350 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15344 17632 16129 17660
rect 15344 17620 15350 17632
rect 16117 17629 16129 17632
rect 16163 17629 16175 17663
rect 16117 17623 16175 17629
rect 10781 17595 10839 17601
rect 9140 17564 9444 17592
rect 5810 17484 5816 17536
rect 5868 17484 5874 17536
rect 6733 17527 6791 17533
rect 6733 17493 6745 17527
rect 6779 17524 6791 17527
rect 7190 17524 7196 17536
rect 6779 17496 7196 17524
rect 6779 17493 6791 17496
rect 6733 17487 6791 17493
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 7834 17524 7840 17536
rect 7524 17496 7840 17524
rect 7524 17484 7530 17496
rect 7834 17484 7840 17496
rect 7892 17484 7898 17536
rect 7926 17484 7932 17536
rect 7984 17484 7990 17536
rect 8386 17484 8392 17536
rect 8444 17524 8450 17536
rect 9140 17533 9168 17564
rect 9125 17527 9183 17533
rect 9125 17524 9137 17527
rect 8444 17496 9137 17524
rect 8444 17484 8450 17496
rect 9125 17493 9137 17496
rect 9171 17493 9183 17527
rect 9125 17487 9183 17493
rect 9306 17484 9312 17536
rect 9364 17484 9370 17536
rect 9416 17524 9444 17564
rect 10781 17561 10793 17595
rect 10827 17561 10839 17595
rect 10781 17555 10839 17561
rect 11057 17527 11115 17533
rect 11057 17524 11069 17527
rect 9416 17496 11069 17524
rect 11057 17493 11069 17496
rect 11103 17493 11115 17527
rect 11057 17487 11115 17493
rect 17862 17484 17868 17536
rect 17920 17484 17926 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 4065 17323 4123 17329
rect 4065 17289 4077 17323
rect 4111 17320 4123 17323
rect 4338 17320 4344 17332
rect 4111 17292 4344 17320
rect 4111 17289 4123 17292
rect 4065 17283 4123 17289
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7098 17320 7104 17332
rect 6963 17292 7104 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 7984 17292 8769 17320
rect 7984 17280 7990 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 8938 17280 8944 17332
rect 8996 17320 9002 17332
rect 11330 17320 11336 17332
rect 8996 17292 11336 17320
rect 8996 17280 9002 17292
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 6089 17255 6147 17261
rect 6089 17221 6101 17255
rect 6135 17252 6147 17255
rect 7006 17252 7012 17264
rect 6135 17224 7012 17252
rect 6135 17221 6147 17224
rect 6089 17215 6147 17221
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 8570 17252 8576 17264
rect 7116 17224 8576 17252
rect 4246 17144 4252 17196
rect 4304 17184 4310 17196
rect 4433 17187 4491 17193
rect 4433 17184 4445 17187
rect 4304 17156 4445 17184
rect 4304 17144 4310 17156
rect 4433 17153 4445 17156
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 5718 17144 5724 17196
rect 5776 17184 5782 17196
rect 7116 17193 7144 17224
rect 8570 17212 8576 17224
rect 8628 17212 8634 17264
rect 10410 17252 10416 17264
rect 9876 17224 10416 17252
rect 7101 17187 7159 17193
rect 5776 17156 6040 17184
rect 5776 17144 5782 17156
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 1912 17088 2329 17116
rect 1912 17076 1918 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 3694 17116 3700 17128
rect 2547 17088 3700 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 3878 17076 3884 17128
rect 3936 17076 3942 17128
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4111 17088 4476 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4448 17057 4476 17088
rect 4614 17076 4620 17128
rect 4672 17076 4678 17128
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17116 4767 17119
rect 5810 17116 5816 17128
rect 4755 17088 5816 17116
rect 4755 17085 4767 17088
rect 4709 17079 4767 17085
rect 5810 17076 5816 17088
rect 5868 17076 5874 17128
rect 6012 17125 6040 17156
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7340 17156 7573 17184
rect 7340 17144 7346 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9493 17187 9551 17193
rect 9493 17184 9505 17187
rect 9364 17156 9505 17184
rect 9364 17144 9370 17156
rect 9493 17153 9505 17156
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9582 17144 9588 17196
rect 9640 17184 9646 17196
rect 9876 17193 9904 17224
rect 10410 17212 10416 17224
rect 10468 17212 10474 17264
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9640 17156 9873 17184
rect 9640 17144 9646 17156
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 10318 17184 10324 17196
rect 9999 17156 10324 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 5997 17079 6055 17085
rect 6270 17076 6276 17128
rect 6328 17076 6334 17128
rect 7193 17119 7251 17125
rect 7193 17085 7205 17119
rect 7239 17116 7251 17119
rect 7374 17116 7380 17128
rect 7239 17088 7380 17116
rect 7239 17085 7251 17088
rect 7193 17079 7251 17085
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9674 17116 9680 17128
rect 8895 17088 9680 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 10134 17076 10140 17128
rect 10192 17076 10198 17128
rect 10229 17119 10287 17125
rect 10229 17085 10241 17119
rect 10275 17085 10287 17119
rect 10229 17079 10287 17085
rect 4433 17051 4491 17057
rect 4433 17017 4445 17051
rect 4479 17017 4491 17051
rect 4433 17011 4491 17017
rect 8662 17008 8668 17060
rect 8720 17048 8726 17060
rect 10244 17048 10272 17079
rect 10410 17076 10416 17128
rect 10468 17076 10474 17128
rect 8720 17020 10272 17048
rect 8720 17008 8726 17020
rect 10686 17008 10692 17060
rect 10744 17048 10750 17060
rect 11241 17051 11299 17057
rect 11241 17048 11253 17051
rect 10744 17020 11253 17048
rect 10744 17008 10750 17020
rect 11241 17017 11253 17020
rect 11287 17048 11299 17051
rect 16758 17048 16764 17060
rect 11287 17020 16764 17048
rect 11287 17017 11299 17020
rect 11241 17011 11299 17017
rect 16758 17008 16764 17020
rect 16816 17048 16822 17060
rect 17862 17048 17868 17060
rect 16816 17020 17868 17048
rect 16816 17008 16822 17020
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 2406 16940 2412 16992
rect 2464 16940 2470 16992
rect 6365 16983 6423 16989
rect 6365 16949 6377 16983
rect 6411 16980 6423 16983
rect 7190 16980 7196 16992
rect 6411 16952 7196 16980
rect 6411 16949 6423 16952
rect 6365 16943 6423 16949
rect 7190 16940 7196 16952
rect 7248 16940 7254 16992
rect 10318 16940 10324 16992
rect 10376 16940 10382 16992
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 4154 16776 4160 16788
rect 2056 16748 4160 16776
rect 2056 16584 2084 16748
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 9674 16776 9680 16788
rect 9539 16748 9680 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 2308 16711 2366 16717
rect 2308 16677 2320 16711
rect 2354 16708 2366 16711
rect 2406 16708 2412 16720
rect 2354 16680 2412 16708
rect 2354 16677 2366 16680
rect 2308 16671 2366 16677
rect 2406 16668 2412 16680
rect 2464 16668 2470 16720
rect 3694 16668 3700 16720
rect 3752 16668 3758 16720
rect 7374 16668 7380 16720
rect 7432 16708 7438 16720
rect 8018 16708 8024 16720
rect 7432 16680 8024 16708
rect 7432 16668 7438 16680
rect 8018 16668 8024 16680
rect 8076 16708 8082 16720
rect 11238 16708 11244 16720
rect 8076 16680 11244 16708
rect 8076 16668 8082 16680
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 3970 16600 3976 16652
rect 4028 16600 4034 16652
rect 4154 16600 4160 16652
rect 4212 16600 4218 16652
rect 4430 16649 4436 16652
rect 4424 16603 4436 16649
rect 4430 16600 4436 16603
rect 4488 16600 4494 16652
rect 9490 16600 9496 16652
rect 9548 16640 9554 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9548 16612 9689 16640
rect 9548 16600 9554 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 10042 16600 10048 16652
rect 10100 16600 10106 16652
rect 2038 16532 2044 16584
rect 2096 16532 2102 16584
rect 3697 16575 3755 16581
rect 3697 16541 3709 16575
rect 3743 16572 3755 16575
rect 5718 16572 5724 16584
rect 3743 16544 4200 16572
rect 3743 16541 3755 16544
rect 3697 16535 3755 16541
rect 4172 16516 4200 16544
rect 5552 16544 5724 16572
rect 3421 16507 3479 16513
rect 3421 16473 3433 16507
rect 3467 16504 3479 16507
rect 3602 16504 3608 16516
rect 3467 16476 3608 16504
rect 3467 16473 3479 16476
rect 3421 16467 3479 16473
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 4154 16464 4160 16516
rect 4212 16464 4218 16516
rect 5552 16513 5580 16544
rect 5718 16532 5724 16544
rect 5776 16572 5782 16584
rect 6365 16575 6423 16581
rect 6365 16572 6377 16575
rect 5776 16544 6377 16572
rect 5776 16532 5782 16544
rect 6365 16541 6377 16544
rect 6411 16541 6423 16575
rect 6365 16535 6423 16541
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16473 5595 16507
rect 5537 16467 5595 16473
rect 3510 16396 3516 16448
rect 3568 16436 3574 16448
rect 3878 16436 3884 16448
rect 3568 16408 3884 16436
rect 3568 16396 3574 16408
rect 3878 16396 3884 16408
rect 3936 16396 3942 16448
rect 5810 16396 5816 16448
rect 5868 16396 5874 16448
rect 7006 16396 7012 16448
rect 7064 16436 7070 16448
rect 8202 16436 8208 16448
rect 7064 16408 8208 16436
rect 7064 16396 7070 16408
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 10686 16436 10692 16448
rect 9999 16408 10692 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 10686 16396 10692 16408
rect 10744 16396 10750 16448
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 3970 16232 3976 16244
rect 3743 16204 3976 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 3970 16192 3976 16204
rect 4028 16192 4034 16244
rect 4709 16235 4767 16241
rect 4709 16201 4721 16235
rect 4755 16232 4767 16235
rect 5442 16232 5448 16244
rect 4755 16204 5448 16232
rect 4755 16201 4767 16204
rect 4709 16195 4767 16201
rect 5442 16192 5448 16204
rect 5500 16192 5506 16244
rect 10042 16232 10048 16244
rect 5828 16204 10048 16232
rect 3510 16124 3516 16176
rect 3568 16164 3574 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 3568 16136 4537 16164
rect 3568 16124 3574 16136
rect 4525 16133 4537 16136
rect 4571 16133 4583 16167
rect 4525 16127 4583 16133
rect 4614 16124 4620 16176
rect 4672 16164 4678 16176
rect 4985 16167 5043 16173
rect 4985 16164 4997 16167
rect 4672 16136 4997 16164
rect 4672 16124 4678 16136
rect 4985 16133 4997 16136
rect 5031 16133 5043 16167
rect 4985 16127 5043 16133
rect 2041 16099 2099 16105
rect 2041 16096 2053 16099
rect 1780 16068 2053 16096
rect 1780 16037 1808 16068
rect 2041 16065 2053 16068
rect 2087 16096 2099 16099
rect 2866 16096 2872 16108
rect 2087 16068 2872 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2866 16056 2872 16068
rect 2924 16056 2930 16108
rect 5442 16096 5448 16108
rect 5184 16068 5448 16096
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 15997 1455 16031
rect 1397 15991 1455 15997
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 1412 15960 1440 15991
rect 1854 15988 1860 16040
rect 1912 15988 1918 16040
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 2832 16000 3433 16028
rect 2832 15988 2838 16000
rect 3421 15997 3433 16000
rect 3467 16028 3479 16031
rect 3510 16028 3516 16040
rect 3467 16000 3516 16028
rect 3467 15997 3479 16000
rect 3421 15991 3479 15997
rect 3510 15988 3516 16000
rect 3568 15988 3574 16040
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 5184 16037 5212 16068
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 5828 16105 5856 16204
rect 10042 16192 10048 16204
rect 10100 16232 10106 16244
rect 10505 16235 10563 16241
rect 10505 16232 10517 16235
rect 10100 16204 10517 16232
rect 10100 16192 10106 16204
rect 10505 16201 10517 16204
rect 10551 16201 10563 16235
rect 10505 16195 10563 16201
rect 11330 16192 11336 16244
rect 11388 16232 11394 16244
rect 12526 16232 12532 16244
rect 11388 16204 12532 16232
rect 11388 16192 11394 16204
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 13170 16192 13176 16244
rect 13228 16192 13234 16244
rect 7926 16124 7932 16176
rect 7984 16124 7990 16176
rect 12434 16124 12440 16176
rect 12492 16164 12498 16176
rect 12621 16167 12679 16173
rect 12621 16164 12633 16167
rect 12492 16136 12633 16164
rect 12492 16124 12498 16136
rect 12621 16133 12633 16136
rect 12667 16164 12679 16167
rect 12667 16136 14412 16164
rect 12667 16133 12679 16136
rect 12621 16127 12679 16133
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 6089 16099 6147 16105
rect 6089 16065 6101 16099
rect 6135 16096 6147 16099
rect 7006 16096 7012 16108
rect 6135 16068 7012 16096
rect 6135 16065 6147 16068
rect 6089 16059 6147 16065
rect 7006 16056 7012 16068
rect 7064 16056 7070 16108
rect 7098 16056 7104 16108
rect 7156 16056 7162 16108
rect 7944 16096 7972 16124
rect 7300 16068 7972 16096
rect 4341 16031 4399 16037
rect 4341 16028 4353 16031
rect 3660 16000 4353 16028
rect 3660 15988 3666 16000
rect 4341 15997 4353 16000
rect 4387 16028 4399 16031
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4387 16000 4660 16028
rect 4387 15997 4399 16000
rect 4341 15991 4399 15997
rect 1872 15960 1900 15988
rect 1412 15932 1808 15960
rect 1872 15932 2774 15960
rect 1670 15852 1676 15904
rect 1728 15852 1734 15904
rect 1780 15892 1808 15932
rect 2314 15892 2320 15904
rect 1780 15864 2320 15892
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 2590 15852 2596 15904
rect 2648 15852 2654 15904
rect 2746 15892 2774 15932
rect 2958 15920 2964 15972
rect 3016 15960 3022 15972
rect 3620 15960 3648 15988
rect 3016 15932 3648 15960
rect 3016 15920 3022 15932
rect 3237 15895 3295 15901
rect 3237 15892 3249 15895
rect 2746 15864 3249 15892
rect 3237 15861 3249 15864
rect 3283 15892 3295 15895
rect 3326 15892 3332 15904
rect 3283 15864 3332 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 3326 15852 3332 15864
rect 3384 15852 3390 15904
rect 4632 15892 4660 16000
rect 4816 16000 5181 16028
rect 4693 15963 4751 15969
rect 4693 15929 4705 15963
rect 4739 15960 4751 15963
rect 4816 15960 4844 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5169 15991 5227 15997
rect 5353 16031 5411 16037
rect 5353 15997 5365 16031
rect 5399 16028 5411 16031
rect 5718 16028 5724 16040
rect 5399 16000 5724 16028
rect 5399 15997 5411 16000
rect 5353 15991 5411 15997
rect 4739 15932 4844 15960
rect 4893 15963 4951 15969
rect 4739 15929 4751 15932
rect 4693 15923 4751 15929
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 5368 15960 5396 15991
rect 5718 15988 5724 16000
rect 5776 15988 5782 16040
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 7213 16031 7271 16037
rect 6512 16000 7144 16028
rect 6512 15988 6518 16000
rect 4939 15932 5396 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 6638 15920 6644 15972
rect 6696 15960 6702 15972
rect 7116 15969 7144 16000
rect 7213 15997 7225 16031
rect 7259 16028 7271 16031
rect 7300 16028 7328 16068
rect 7259 16000 7328 16028
rect 7259 15997 7271 16000
rect 7213 15991 7271 15997
rect 7374 15988 7380 16040
rect 7432 15988 7438 16040
rect 7576 16037 7604 16068
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13136 16068 13553 16096
rect 13136 16056 13142 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 14384 16040 14412 16136
rect 7561 16031 7619 16037
rect 7561 15997 7573 16031
rect 7607 15997 7619 16031
rect 7561 15991 7619 15997
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 15997 7711 16031
rect 7653 15991 7711 15997
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 7929 16031 7987 16037
rect 7929 15997 7941 16031
rect 7975 16028 7987 16031
rect 8110 16028 8116 16040
rect 7975 16000 8116 16028
rect 7975 15997 7987 16000
rect 7929 15991 7987 15997
rect 6825 15963 6883 15969
rect 6825 15960 6837 15963
rect 6696 15932 6837 15960
rect 6696 15920 6702 15932
rect 6825 15929 6837 15932
rect 6871 15929 6883 15963
rect 6825 15923 6883 15929
rect 7009 15963 7067 15969
rect 7009 15929 7021 15963
rect 7055 15929 7067 15963
rect 7009 15923 7067 15929
rect 7101 15963 7159 15969
rect 7101 15929 7113 15963
rect 7147 15960 7159 15963
rect 7668 15960 7696 15991
rect 7147 15932 7696 15960
rect 7760 15960 7788 15991
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 9122 15988 9128 16040
rect 9180 15988 9186 16040
rect 11054 15988 11060 16040
rect 11112 15988 11118 16040
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 13817 16031 13875 16037
rect 13817 16028 13829 16031
rect 13320 16000 13829 16028
rect 13320 15988 13326 16000
rect 13817 15997 13829 16000
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14366 15988 14372 16040
rect 14424 15988 14430 16040
rect 14553 16031 14611 16037
rect 14553 15997 14565 16031
rect 14599 16028 14611 16031
rect 14918 16028 14924 16040
rect 14599 16000 14924 16028
rect 14599 15997 14611 16000
rect 14553 15991 14611 15997
rect 14918 15988 14924 16000
rect 14976 15988 14982 16040
rect 8386 15960 8392 15972
rect 7760 15932 8392 15960
rect 7147 15929 7159 15932
rect 7101 15923 7159 15929
rect 6656 15892 6684 15920
rect 4632 15864 6684 15892
rect 7024 15892 7052 15923
rect 8386 15920 8392 15932
rect 8444 15920 8450 15972
rect 9214 15920 9220 15972
rect 9272 15960 9278 15972
rect 9370 15963 9428 15969
rect 9370 15960 9382 15963
rect 9272 15932 9382 15960
rect 9272 15920 9278 15932
rect 9370 15929 9382 15932
rect 9416 15929 9428 15963
rect 9370 15923 9428 15929
rect 12894 15920 12900 15972
rect 12952 15960 12958 15972
rect 12989 15963 13047 15969
rect 12989 15960 13001 15963
rect 12952 15932 13001 15960
rect 12952 15920 12958 15932
rect 12989 15929 13001 15932
rect 13035 15929 13047 15963
rect 12989 15923 13047 15929
rect 13446 15920 13452 15972
rect 13504 15960 13510 15972
rect 13909 15963 13967 15969
rect 13909 15960 13921 15963
rect 13504 15932 13921 15960
rect 13504 15920 13510 15932
rect 13909 15929 13921 15932
rect 13955 15960 13967 15963
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 13955 15932 14197 15960
rect 13955 15929 13967 15932
rect 13909 15923 13967 15929
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 14185 15923 14243 15929
rect 7190 15892 7196 15904
rect 7024 15864 7196 15892
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 8113 15895 8171 15901
rect 8113 15861 8125 15895
rect 8159 15892 8171 15895
rect 11974 15892 11980 15904
rect 8159 15864 11980 15892
rect 8159 15861 8171 15864
rect 8113 15855 8171 15861
rect 11974 15852 11980 15864
rect 12032 15892 12038 15904
rect 12342 15892 12348 15904
rect 12032 15864 12348 15892
rect 12032 15852 12038 15864
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13189 15895 13247 15901
rect 13189 15892 13201 15895
rect 12860 15864 13201 15892
rect 12860 15852 12866 15864
rect 13189 15861 13201 15864
rect 13235 15861 13247 15895
rect 13189 15855 13247 15861
rect 13354 15852 13360 15904
rect 13412 15852 13418 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13596 15864 13737 15892
rect 13596 15852 13602 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 14090 15852 14096 15904
rect 14148 15852 14154 15904
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 3697 15691 3755 15697
rect 3697 15688 3709 15691
rect 1596 15660 3709 15688
rect 1596 15552 1624 15660
rect 3697 15657 3709 15660
rect 3743 15657 3755 15691
rect 3697 15651 3755 15657
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4617 15691 4675 15697
rect 4617 15688 4629 15691
rect 4488 15660 4629 15688
rect 4488 15648 4494 15660
rect 4617 15657 4629 15660
rect 4663 15657 4675 15691
rect 4617 15651 4675 15657
rect 6914 15648 6920 15700
rect 6972 15648 6978 15700
rect 7193 15691 7251 15697
rect 7193 15657 7205 15691
rect 7239 15688 7251 15691
rect 7374 15688 7380 15700
rect 7239 15660 7380 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7524 15660 7573 15688
rect 7524 15648 7530 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 7561 15651 7619 15657
rect 9214 15648 9220 15700
rect 9272 15648 9278 15700
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 9861 15691 9919 15697
rect 9861 15688 9873 15691
rect 9732 15660 9873 15688
rect 9732 15648 9738 15660
rect 9861 15657 9873 15660
rect 9907 15657 9919 15691
rect 9861 15651 9919 15657
rect 11330 15648 11336 15700
rect 11388 15648 11394 15700
rect 12802 15648 12808 15700
rect 12860 15648 12866 15700
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 15286 15688 15292 15700
rect 13688 15660 15292 15688
rect 13688 15648 13694 15660
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 1670 15580 1676 15632
rect 1728 15620 1734 15632
rect 4157 15623 4215 15629
rect 1728 15592 3556 15620
rect 1728 15580 1734 15592
rect 1958 15555 2016 15561
rect 1958 15552 1970 15555
rect 1596 15524 1970 15552
rect 1958 15521 1970 15524
rect 2004 15521 2016 15555
rect 1958 15515 2016 15521
rect 2130 15512 2136 15564
rect 2188 15552 2194 15564
rect 2225 15555 2283 15561
rect 2225 15552 2237 15555
rect 2188 15524 2237 15552
rect 2188 15512 2194 15524
rect 2225 15521 2237 15524
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2590 15512 2596 15564
rect 2648 15552 2654 15564
rect 3237 15555 3295 15561
rect 3237 15552 3249 15555
rect 2648 15524 3249 15552
rect 2648 15512 2654 15524
rect 3237 15521 3249 15524
rect 3283 15521 3295 15555
rect 3237 15515 3295 15521
rect 3326 15512 3332 15564
rect 3384 15512 3390 15564
rect 3528 15561 3556 15592
rect 4157 15589 4169 15623
rect 4203 15620 4215 15623
rect 6932 15620 6960 15648
rect 4203 15592 4568 15620
rect 6932 15592 7052 15620
rect 4203 15589 4215 15592
rect 4157 15583 4215 15589
rect 4540 15561 4568 15592
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15521 3571 15555
rect 3513 15515 3571 15521
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 2774 15444 2780 15496
rect 2832 15444 2838 15496
rect 2866 15444 2872 15496
rect 2924 15444 2930 15496
rect 2958 15444 2964 15496
rect 3016 15444 3022 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3142 15484 3148 15496
rect 3099 15456 3148 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4448 15484 4476 15515
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4672 15524 4721 15552
rect 4672 15512 4678 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 6730 15552 6736 15564
rect 6687 15524 6736 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 7024 15561 7052 15592
rect 7282 15580 7288 15632
rect 7340 15620 7346 15632
rect 11698 15620 11704 15632
rect 7340 15592 11704 15620
rect 7340 15580 7346 15592
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 11808 15592 12756 15620
rect 11808 15564 11836 15592
rect 6917 15555 6975 15561
rect 6917 15521 6929 15555
rect 6963 15521 6975 15555
rect 6917 15515 6975 15521
rect 7009 15555 7067 15561
rect 7009 15521 7021 15555
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 5810 15484 5816 15496
rect 4448 15456 5816 15484
rect 5810 15444 5816 15456
rect 5868 15444 5874 15496
rect 6932 15484 6960 15515
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7444 15555 7502 15561
rect 7444 15552 7456 15555
rect 7156 15524 7456 15552
rect 7156 15512 7162 15524
rect 7444 15521 7456 15524
rect 7490 15521 7502 15555
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7444 15515 7502 15521
rect 7576 15524 8033 15552
rect 7576 15484 7604 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8202 15512 8208 15564
rect 8260 15512 8266 15564
rect 8294 15512 8300 15564
rect 8352 15512 8358 15564
rect 8386 15512 8392 15564
rect 8444 15512 8450 15564
rect 8665 15555 8723 15561
rect 8665 15521 8677 15555
rect 8711 15552 8723 15555
rect 8938 15552 8944 15564
rect 8711 15524 8944 15552
rect 8711 15521 8723 15524
rect 8665 15515 8723 15521
rect 8938 15512 8944 15524
rect 8996 15512 9002 15564
rect 9398 15512 9404 15564
rect 9456 15512 9462 15564
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15552 9551 15555
rect 9582 15552 9588 15564
rect 9539 15524 9588 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 9582 15512 9588 15524
rect 9640 15512 9646 15564
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 5920 15456 7604 15484
rect 7653 15487 7711 15493
rect 2884 15416 2912 15444
rect 3234 15416 3240 15428
rect 2332 15388 3240 15416
rect 845 15351 903 15357
rect 845 15317 857 15351
rect 891 15348 903 15351
rect 2332 15348 2360 15388
rect 3234 15376 3240 15388
rect 3292 15416 3298 15428
rect 5920 15416 5948 15456
rect 7653 15453 7665 15487
rect 7699 15484 7711 15487
rect 7834 15484 7840 15496
rect 7699 15456 7840 15484
rect 7699 15453 7711 15456
rect 7653 15447 7711 15453
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15453 8815 15487
rect 8757 15447 8815 15453
rect 3292 15388 5948 15416
rect 6733 15419 6791 15425
rect 3292 15376 3298 15388
rect 6733 15385 6745 15419
rect 6779 15416 6791 15419
rect 7944 15416 7972 15447
rect 8573 15419 8631 15425
rect 8573 15416 8585 15419
rect 6779 15388 7880 15416
rect 7944 15388 8585 15416
rect 6779 15385 6791 15388
rect 6733 15379 6791 15385
rect 891 15320 2360 15348
rect 891 15317 903 15320
rect 845 15311 903 15317
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 2593 15351 2651 15357
rect 2593 15348 2605 15351
rect 2464 15320 2605 15348
rect 2464 15308 2470 15320
rect 2593 15317 2605 15320
rect 2639 15317 2651 15351
rect 2593 15311 2651 15317
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 5442 15348 5448 15360
rect 4387 15320 5448 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 7282 15308 7288 15360
rect 7340 15308 7346 15360
rect 7852 15348 7880 15388
rect 8573 15385 8585 15388
rect 8619 15385 8631 15419
rect 8772 15416 8800 15447
rect 9490 15416 9496 15428
rect 8772 15388 9496 15416
rect 8573 15379 8631 15385
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 8018 15348 8024 15360
rect 7852 15320 8024 15348
rect 8018 15308 8024 15320
rect 8076 15348 8082 15360
rect 8665 15351 8723 15357
rect 8665 15348 8677 15351
rect 8076 15320 8677 15348
rect 8076 15308 8082 15320
rect 8665 15317 8677 15320
rect 8711 15317 8723 15351
rect 8665 15311 8723 15317
rect 9030 15308 9036 15360
rect 9088 15308 9094 15360
rect 11532 15348 11560 15515
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12434 15552 12440 15564
rect 12023 15524 12440 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 12526 15512 12532 15564
rect 12584 15512 12590 15564
rect 12728 15561 12756 15592
rect 13354 15580 13360 15632
rect 13412 15620 13418 15632
rect 13412 15592 15240 15620
rect 13412 15580 13418 15592
rect 12713 15555 12771 15561
rect 12713 15521 12725 15555
rect 12759 15521 12771 15555
rect 12713 15515 12771 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13004 15552 13124 15556
rect 12943 15528 13400 15552
rect 12943 15524 13032 15528
rect 13096 15524 13400 15528
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 12084 15456 12265 15484
rect 11698 15376 11704 15428
rect 11756 15416 11762 15428
rect 12084 15416 12112 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 11756 15388 12112 15416
rect 11756 15376 11762 15388
rect 12069 15351 12127 15357
rect 12069 15348 12081 15351
rect 11532 15320 12081 15348
rect 12069 15317 12081 15320
rect 12115 15317 12127 15351
rect 12069 15311 12127 15317
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 13188 15348 13216 15447
rect 13262 15444 13268 15496
rect 13320 15444 13326 15496
rect 13372 15493 13400 15524
rect 13630 15512 13636 15564
rect 13688 15512 13694 15564
rect 13906 15561 13912 15564
rect 13900 15515 13912 15561
rect 13906 15512 13912 15515
rect 13964 15512 13970 15564
rect 15212 15561 15240 15592
rect 15197 15555 15255 15561
rect 15197 15521 15209 15555
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13446 15484 13452 15496
rect 13403 15456 13452 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 13446 15348 13452 15360
rect 13136 15320 13452 15348
rect 13136 15308 13142 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13630 15348 13636 15360
rect 13587 15320 13636 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 15102 15348 15108 15360
rect 15059 15320 15108 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15378 15308 15384 15360
rect 15436 15308 15442 15360
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 2314 15104 2320 15156
rect 2372 15144 2378 15156
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 2372 15116 2421 15144
rect 2372 15104 2378 15116
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 2409 15107 2467 15113
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3142 15144 3148 15156
rect 2915 15116 3148 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3142 15104 3148 15116
rect 3200 15144 3206 15156
rect 3510 15144 3516 15156
rect 3200 15116 3516 15144
rect 3200 15104 3206 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 6178 15104 6184 15156
rect 6236 15144 6242 15156
rect 11149 15147 11207 15153
rect 11149 15144 11161 15147
rect 6236 15116 11161 15144
rect 6236 15104 6242 15116
rect 11149 15113 11161 15116
rect 11195 15113 11207 15147
rect 11149 15107 11207 15113
rect 11517 15147 11575 15153
rect 11517 15113 11529 15147
rect 11563 15144 11575 15147
rect 11790 15144 11796 15156
rect 11563 15116 11796 15144
rect 11563 15113 11575 15116
rect 11517 15107 11575 15113
rect 1670 15036 1676 15088
rect 1728 15076 1734 15088
rect 2041 15079 2099 15085
rect 2041 15076 2053 15079
rect 1728 15048 2053 15076
rect 1728 15036 1734 15048
rect 2041 15045 2053 15048
rect 2087 15076 2099 15079
rect 2685 15079 2743 15085
rect 2685 15076 2697 15079
rect 2087 15048 2697 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 2685 15045 2697 15048
rect 2731 15045 2743 15079
rect 2685 15039 2743 15045
rect 2314 14968 2320 15020
rect 2372 15008 2378 15020
rect 4154 15008 4160 15020
rect 2372 14980 4160 15008
rect 2372 14968 2378 14980
rect 4154 14968 4160 14980
rect 4212 15008 4218 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4212 14980 4905 15008
rect 4212 14968 4218 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 6362 14900 6368 14952
rect 6420 14940 6426 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 6420 14912 6653 14940
rect 6420 14900 6426 14912
rect 6641 14909 6653 14912
rect 6687 14940 6699 14943
rect 9122 14940 9128 14952
rect 6687 14912 9128 14940
rect 6687 14909 6699 14912
rect 6641 14903 6699 14909
rect 9122 14900 9128 14912
rect 9180 14940 9186 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9180 14912 9965 14940
rect 9180 14900 9186 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 10686 14900 10692 14952
rect 10744 14940 10750 14952
rect 10965 14943 11023 14949
rect 10965 14940 10977 14943
rect 10744 14912 10977 14940
rect 10744 14900 10750 14912
rect 10965 14909 10977 14912
rect 11011 14909 11023 14943
rect 10965 14903 11023 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 11532 14940 11560 15107
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 12805 15147 12863 15153
rect 12805 15113 12817 15147
rect 12851 15144 12863 15147
rect 13170 15144 13176 15156
rect 12851 15116 13176 15144
rect 12851 15113 12863 15116
rect 12805 15107 12863 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 14918 15144 14924 15156
rect 13372 15116 14924 15144
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 11974 15008 11980 15020
rect 11931 14980 11980 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 11974 14968 11980 14980
rect 12032 15008 12038 15020
rect 13078 15008 13084 15020
rect 12032 14980 13084 15008
rect 12032 14968 12038 14980
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 13372 15008 13400 15116
rect 14918 15104 14924 15116
rect 14976 15104 14982 15156
rect 15102 15104 15108 15156
rect 15160 15144 15166 15156
rect 16850 15144 16856 15156
rect 15160 15116 16856 15144
rect 15160 15104 15166 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 14139 15079 14197 15085
rect 14139 15076 14151 15079
rect 13504 15048 14151 15076
rect 13504 15036 13510 15048
rect 14139 15045 14151 15048
rect 14185 15045 14197 15079
rect 14139 15039 14197 15045
rect 14458 15036 14464 15088
rect 14516 15076 14522 15088
rect 15120 15076 15148 15104
rect 14516 15048 15148 15076
rect 14516 15036 14522 15048
rect 15105 15011 15163 15017
rect 13311 14980 13400 15008
rect 13464 14980 13860 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 11195 14912 11560 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 12986 14940 12992 14952
rect 11756 14912 12992 14940
rect 11756 14900 11762 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 13173 14943 13231 14949
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 13464 14940 13492 14980
rect 13219 14912 13492 14940
rect 13541 14943 13599 14949
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13541 14903 13599 14909
rect 2406 14832 2412 14884
rect 2464 14832 2470 14884
rect 3053 14875 3111 14881
rect 3053 14841 3065 14875
rect 3099 14872 3111 14875
rect 3234 14872 3240 14884
rect 3099 14844 3240 14872
rect 3099 14841 3111 14844
rect 3053 14835 3111 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 5077 14875 5135 14881
rect 5077 14841 5089 14875
rect 5123 14872 5135 14875
rect 6178 14872 6184 14884
rect 5123 14844 6184 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 6178 14832 6184 14844
rect 6236 14832 6242 14884
rect 7098 14832 7104 14884
rect 7156 14872 7162 14884
rect 8205 14875 8263 14881
rect 8205 14872 8217 14875
rect 7156 14844 8217 14872
rect 7156 14832 7162 14844
rect 8205 14841 8217 14844
rect 8251 14841 8263 14875
rect 8205 14835 8263 14841
rect 9490 14832 9496 14884
rect 9548 14872 9554 14884
rect 9686 14875 9744 14881
rect 9686 14872 9698 14875
rect 9548 14844 9698 14872
rect 9548 14832 9554 14844
rect 9686 14841 9698 14844
rect 9732 14841 9744 14875
rect 9686 14835 9744 14841
rect 10781 14875 10839 14881
rect 10781 14841 10793 14875
rect 10827 14872 10839 14875
rect 11514 14872 11520 14884
rect 10827 14844 11520 14872
rect 10827 14841 10839 14844
rect 10781 14835 10839 14841
rect 11514 14832 11520 14844
rect 11572 14872 11578 14884
rect 12894 14872 12900 14884
rect 11572 14844 12900 14872
rect 11572 14832 11578 14844
rect 12894 14832 12900 14844
rect 12952 14872 12958 14884
rect 13556 14872 13584 14903
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 13688 14912 13737 14940
rect 13688 14900 13694 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 12952 14844 13584 14872
rect 13832 14872 13860 14980
rect 15105 14977 15117 15011
rect 15151 15008 15163 15011
rect 15286 15008 15292 15020
rect 15151 14980 15292 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15378 14968 15384 15020
rect 15436 14968 15442 15020
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 14090 14940 14096 14952
rect 13955 14912 14096 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 14090 14900 14096 14912
rect 14148 14900 14154 14952
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 16816 14912 16865 14940
rect 16816 14900 16822 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 16942 14900 16948 14952
rect 17000 14900 17006 14952
rect 14366 14872 14372 14884
rect 13832 14844 14372 14872
rect 12952 14832 12958 14844
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 17402 14872 17408 14884
rect 16684 14844 17408 14872
rect 2130 14764 2136 14816
rect 2188 14804 2194 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 2188 14776 2605 14804
rect 2188 14764 2194 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2593 14767 2651 14773
rect 2853 14807 2911 14813
rect 2853 14773 2865 14807
rect 2899 14804 2911 14807
rect 3326 14804 3332 14816
rect 2899 14776 3332 14804
rect 2899 14773 2911 14776
rect 2853 14767 2911 14773
rect 3326 14764 3332 14776
rect 3384 14764 3390 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8573 14807 8631 14813
rect 8573 14804 8585 14807
rect 8168 14776 8585 14804
rect 8168 14764 8174 14776
rect 8573 14773 8585 14776
rect 8619 14773 8631 14807
rect 8573 14767 8631 14773
rect 13538 14764 13544 14816
rect 13596 14764 13602 14816
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 16684 14813 16712 14844
rect 17402 14832 17408 14844
rect 17460 14832 17466 14884
rect 16669 14807 16727 14813
rect 16669 14804 16681 14807
rect 14976 14776 16681 14804
rect 14976 14764 14982 14776
rect 16669 14773 16681 14776
rect 16715 14773 16727 14807
rect 16669 14767 16727 14773
rect 17126 14764 17132 14816
rect 17184 14804 17190 14816
rect 17221 14807 17279 14813
rect 17221 14804 17233 14807
rect 17184 14776 17233 14804
rect 17184 14764 17190 14776
rect 17221 14773 17233 14776
rect 17267 14773 17279 14807
rect 17221 14767 17279 14773
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 6825 14603 6883 14609
rect 6825 14600 6837 14603
rect 4172 14572 6837 14600
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2038 14464 2044 14476
rect 1995 14436 2044 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2222 14473 2228 14476
rect 2216 14427 2228 14473
rect 2222 14424 2228 14427
rect 2280 14424 2286 14476
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14464 4031 14467
rect 4062 14464 4068 14476
rect 4019 14436 4068 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4172 14473 4200 14572
rect 6825 14569 6837 14572
rect 6871 14600 6883 14603
rect 7745 14603 7803 14609
rect 6871 14572 7604 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 4709 14535 4767 14541
rect 4709 14501 4721 14535
rect 4755 14532 4767 14535
rect 6178 14532 6184 14544
rect 4755 14504 6184 14532
rect 4755 14501 4767 14504
rect 4709 14495 4767 14501
rect 6178 14492 6184 14504
rect 6236 14492 6242 14544
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14464 4215 14467
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 4203 14436 4261 14464
rect 4203 14433 4215 14436
rect 4157 14427 4215 14433
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4430 14424 4436 14476
rect 4488 14424 4494 14476
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 5169 14427 5227 14433
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14464 5411 14467
rect 5626 14464 5632 14476
rect 5399 14436 5632 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4387 14368 5089 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 5077 14365 5089 14368
rect 5123 14396 5135 14399
rect 5184 14396 5212 14427
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6380 14436 6469 14464
rect 5123 14368 5212 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 4065 14331 4123 14337
rect 4065 14297 4077 14331
rect 4111 14328 4123 14331
rect 4111 14300 4752 14328
rect 4111 14297 4123 14300
rect 4065 14291 4123 14297
rect 3329 14263 3387 14269
rect 3329 14229 3341 14263
rect 3375 14260 3387 14263
rect 3510 14260 3516 14272
rect 3375 14232 3516 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 4525 14263 4583 14269
rect 4525 14229 4537 14263
rect 4571 14260 4583 14263
rect 4614 14260 4620 14272
rect 4571 14232 4620 14260
rect 4571 14229 4583 14232
rect 4525 14223 4583 14229
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 4724 14269 4752 14300
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 6380 14337 6408 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6730 14424 6736 14476
rect 6788 14424 6794 14476
rect 6822 14424 6828 14476
rect 6880 14464 6886 14476
rect 7009 14467 7067 14473
rect 7009 14464 7021 14467
rect 6880 14436 7021 14464
rect 6880 14424 6886 14436
rect 7009 14433 7021 14436
rect 7055 14433 7067 14467
rect 7009 14427 7067 14433
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 7576 14473 7604 14572
rect 7745 14569 7757 14603
rect 7791 14600 7803 14603
rect 7834 14600 7840 14612
rect 7791 14572 7840 14600
rect 7791 14569 7803 14572
rect 7745 14563 7803 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 8018 14560 8024 14612
rect 8076 14560 8082 14612
rect 8849 14603 8907 14609
rect 8849 14569 8861 14603
rect 8895 14600 8907 14603
rect 9030 14600 9036 14612
rect 8895 14572 9036 14600
rect 8895 14569 8907 14572
rect 8849 14563 8907 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9490 14560 9496 14612
rect 9548 14560 9554 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 13906 14600 13912 14612
rect 13495 14572 13912 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 13906 14560 13912 14572
rect 13964 14560 13970 14612
rect 16761 14603 16819 14609
rect 16761 14569 16773 14603
rect 16807 14600 16819 14603
rect 16942 14600 16948 14612
rect 16807 14572 16948 14600
rect 16807 14569 16819 14572
rect 16761 14563 16819 14569
rect 12618 14532 12624 14544
rect 10980 14504 12624 14532
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14433 7619 14467
rect 7561 14427 7619 14433
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 9306 14424 9312 14476
rect 9364 14464 9370 14476
rect 10980 14464 11008 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 16776 14532 16804 14563
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 15028 14504 16804 14532
rect 9364 14436 11008 14464
rect 9364 14424 9370 14436
rect 11146 14424 11152 14476
rect 11204 14464 11210 14476
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11204 14436 11529 14464
rect 11204 14424 11210 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 13357 14467 13415 14473
rect 13357 14433 13369 14467
rect 13403 14464 13415 14467
rect 13446 14464 13452 14476
rect 13403 14436 13452 14464
rect 13403 14433 13415 14436
rect 13357 14427 13415 14433
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 13538 14424 13544 14476
rect 13596 14424 13602 14476
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 15028 14473 15056 14504
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14976 14436 15025 14464
rect 14976 14424 14982 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 15102 14424 15108 14476
rect 15160 14464 15166 14476
rect 15289 14467 15347 14473
rect 15289 14464 15301 14467
rect 15160 14436 15301 14464
rect 15160 14424 15166 14436
rect 15289 14433 15301 14436
rect 15335 14433 15347 14467
rect 15289 14427 15347 14433
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6696 14368 7297 14396
rect 6696 14356 6702 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14396 7435 14399
rect 8128 14396 8156 14424
rect 7423 14368 8156 14396
rect 7423 14365 7435 14368
rect 7377 14359 7435 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8536 14368 9229 14396
rect 8536 14356 8542 14368
rect 9217 14365 9229 14368
rect 9263 14396 9275 14399
rect 9582 14396 9588 14408
rect 9263 14368 9588 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 10836 14368 11253 14396
rect 10836 14356 10842 14368
rect 11241 14365 11253 14368
rect 11287 14396 11299 14399
rect 11287 14368 11560 14396
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 5813 14331 5871 14337
rect 5813 14328 5825 14331
rect 5500 14300 5825 14328
rect 5500 14288 5506 14300
rect 5813 14297 5825 14300
rect 5859 14297 5871 14331
rect 5813 14291 5871 14297
rect 6365 14331 6423 14337
rect 6365 14297 6377 14331
rect 6411 14297 6423 14331
rect 6365 14291 6423 14297
rect 11422 14288 11428 14340
rect 11480 14288 11486 14340
rect 11532 14328 11560 14368
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12161 14399 12219 14405
rect 12161 14396 12173 14399
rect 12124 14368 12173 14396
rect 12124 14356 12130 14368
rect 12161 14365 12173 14368
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14424 14368 15608 14396
rect 14424 14356 14430 14368
rect 14734 14328 14740 14340
rect 11532 14300 14740 14328
rect 14734 14288 14740 14300
rect 14792 14288 14798 14340
rect 4709 14263 4767 14269
rect 4709 14229 4721 14263
rect 4755 14229 4767 14263
rect 4709 14223 4767 14229
rect 5537 14263 5595 14269
rect 5537 14229 5549 14263
rect 5583 14260 5595 14263
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5583 14232 6193 14260
rect 5583 14229 5595 14232
rect 5537 14223 5595 14229
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 6638 14220 6644 14272
rect 6696 14220 6702 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 11296 14232 11345 14260
rect 11296 14220 11302 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 11606 14220 11612 14272
rect 11664 14220 11670 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 13504 14232 15117 14260
rect 13504 14220 13510 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15105 14223 15163 14229
rect 15470 14220 15476 14272
rect 15528 14220 15534 14272
rect 15580 14260 15608 14368
rect 16408 14328 16436 14504
rect 16485 14467 16543 14473
rect 16485 14433 16497 14467
rect 16531 14464 16543 14467
rect 16574 14464 16580 14476
rect 16531 14436 16580 14464
rect 16531 14433 16543 14436
rect 16485 14427 16543 14433
rect 16574 14424 16580 14436
rect 16632 14424 16638 14476
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 16724 14436 16957 14464
rect 16724 14424 16730 14436
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17126 14424 17132 14476
rect 17184 14424 17190 14476
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17402 14464 17408 14476
rect 17267 14436 17408 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 16482 14328 16488 14340
rect 16408 14300 16488 14328
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 17221 14263 17279 14269
rect 17221 14260 17233 14263
rect 15580 14232 17233 14260
rect 17221 14229 17233 14232
rect 17267 14260 17279 14263
rect 17310 14260 17316 14272
rect 17267 14232 17316 14260
rect 17267 14229 17279 14232
rect 17221 14223 17279 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17405 14263 17463 14269
rect 17405 14229 17417 14263
rect 17451 14260 17463 14263
rect 18138 14260 18144 14272
rect 17451 14232 18144 14260
rect 17451 14229 17463 14232
rect 17405 14223 17463 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 2041 14059 2099 14065
rect 2041 14025 2053 14059
rect 2087 14056 2099 14059
rect 2222 14056 2228 14068
rect 2087 14028 2228 14056
rect 2087 14025 2099 14028
rect 2041 14019 2099 14025
rect 2222 14016 2228 14028
rect 2280 14016 2286 14068
rect 5442 14016 5448 14068
rect 5500 14016 5506 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 5684 14028 7757 14056
rect 5684 14016 5690 14028
rect 7745 14025 7757 14028
rect 7791 14056 7803 14059
rect 8202 14056 8208 14068
rect 7791 14028 8208 14056
rect 7791 14025 7803 14028
rect 7745 14019 7803 14025
rect 8202 14016 8208 14028
rect 8260 14016 8266 14068
rect 11422 14016 11428 14068
rect 11480 14056 11486 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 11480 14028 13553 14056
rect 11480 14016 11486 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 13541 14019 13599 14025
rect 15102 14016 15108 14068
rect 15160 14016 15166 14068
rect 16574 14016 16580 14068
rect 16632 14016 16638 14068
rect 2409 13991 2467 13997
rect 2409 13957 2421 13991
rect 2455 13957 2467 13991
rect 2409 13951 2467 13957
rect 5353 13991 5411 13997
rect 5353 13957 5365 13991
rect 5399 13988 5411 13991
rect 17678 13988 17684 14000
rect 5399 13960 5764 13988
rect 5399 13957 5411 13960
rect 5353 13951 5411 13957
rect 2314 13880 2320 13932
rect 2372 13880 2378 13932
rect 2424 13920 2452 13951
rect 2424 13892 2728 13920
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2188 13824 2237 13852
rect 2188 13812 2194 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 2498 13812 2504 13864
rect 2556 13812 2562 13864
rect 2700 13861 2728 13892
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13821 2743 13855
rect 2685 13815 2743 13821
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 3418 13852 3424 13864
rect 2915 13824 3424 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 2608 13784 2636 13815
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 3970 13812 3976 13864
rect 4028 13812 4034 13864
rect 5626 13812 5632 13864
rect 5684 13812 5690 13864
rect 5736 13861 5764 13960
rect 16776 13960 17684 13988
rect 6362 13880 6368 13932
rect 6420 13880 6426 13932
rect 13906 13920 13912 13932
rect 12544 13892 13912 13920
rect 6638 13861 6644 13864
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6632 13852 6644 13861
rect 5767 13824 6132 13852
rect 6599 13824 6644 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 2958 13784 2964 13796
rect 2608 13756 2964 13784
rect 2958 13744 2964 13756
rect 3016 13744 3022 13796
rect 4240 13787 4298 13793
rect 4240 13753 4252 13787
rect 4286 13784 4298 13787
rect 4430 13784 4436 13796
rect 4286 13756 4436 13784
rect 4286 13753 4298 13756
rect 4240 13747 4298 13753
rect 4430 13744 4436 13756
rect 4488 13744 4494 13796
rect 5994 13744 6000 13796
rect 6052 13744 6058 13796
rect 6104 13784 6132 13824
rect 6632 13815 6644 13824
rect 6638 13812 6644 13815
rect 6696 13812 6702 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11149 13855 11207 13861
rect 11149 13852 11161 13855
rect 11112 13824 11161 13852
rect 11112 13812 11118 13824
rect 11149 13821 11161 13824
rect 11195 13821 11207 13855
rect 11149 13815 11207 13821
rect 6730 13784 6736 13796
rect 6104 13756 6736 13784
rect 6730 13744 6736 13756
rect 6788 13744 6794 13796
rect 11164 13784 11192 13815
rect 11238 13812 11244 13864
rect 11296 13852 11302 13864
rect 11405 13855 11463 13861
rect 11405 13852 11417 13855
rect 11296 13824 11417 13852
rect 11296 13812 11302 13824
rect 11405 13821 11417 13824
rect 11451 13821 11463 13855
rect 11405 13815 11463 13821
rect 12544 13784 12572 13892
rect 13906 13880 13912 13892
rect 13964 13920 13970 13932
rect 16776 13929 16804 13960
rect 17678 13948 17684 13960
rect 17736 13948 17742 14000
rect 16761 13923 16819 13929
rect 13964 13892 15240 13920
rect 13964 13880 13970 13892
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 11164 13756 12572 13784
rect 12636 13824 12725 13852
rect 12636 13728 12664 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12713 13815 12771 13821
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 13403 13824 13553 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13541 13815 13599 13821
rect 13740 13824 13829 13852
rect 13446 13784 13452 13796
rect 12728 13756 13452 13784
rect 12728 13728 12756 13756
rect 13446 13744 13452 13756
rect 13504 13784 13510 13796
rect 13740 13784 13768 13824
rect 13817 13821 13829 13824
rect 13863 13852 13875 13855
rect 14829 13855 14887 13861
rect 14829 13852 14841 13855
rect 13863 13824 14841 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 14829 13821 14841 13824
rect 14875 13821 14887 13855
rect 14829 13815 14887 13821
rect 14918 13812 14924 13864
rect 14976 13812 14982 13864
rect 15212 13861 15240 13892
rect 16761 13889 16773 13923
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 17494 13880 17500 13932
rect 17552 13880 17558 13932
rect 15197 13855 15255 13861
rect 15197 13821 15209 13855
rect 15243 13852 15255 13855
rect 15286 13852 15292 13864
rect 15243 13824 15292 13852
rect 15243 13821 15255 13824
rect 15197 13815 15255 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15470 13861 15476 13864
rect 15464 13852 15476 13861
rect 15431 13824 15476 13852
rect 15464 13815 15476 13824
rect 15470 13812 15476 13815
rect 15528 13812 15534 13864
rect 16942 13812 16948 13864
rect 17000 13852 17006 13864
rect 17000 13824 17066 13852
rect 17000 13812 17006 13824
rect 13504 13756 13768 13784
rect 13504 13744 13510 13756
rect 14734 13744 14740 13796
rect 14792 13784 14798 13796
rect 15102 13784 15108 13796
rect 14792 13756 15108 13784
rect 14792 13744 14798 13756
rect 15102 13744 15108 13756
rect 15160 13744 15166 13796
rect 2777 13719 2835 13725
rect 2777 13685 2789 13719
rect 2823 13716 2835 13719
rect 3142 13716 3148 13728
rect 2823 13688 3148 13716
rect 2823 13685 2835 13688
rect 2777 13679 2835 13685
rect 3142 13676 3148 13688
rect 3200 13676 3206 13728
rect 5810 13676 5816 13728
rect 5868 13676 5874 13728
rect 12529 13719 12587 13725
rect 12529 13685 12541 13719
rect 12575 13716 12587 13719
rect 12618 13716 12624 13728
rect 12575 13688 12624 13716
rect 12575 13685 12587 13688
rect 12529 13679 12587 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12710 13676 12716 13728
rect 12768 13676 12774 13728
rect 13722 13676 13728 13728
rect 13780 13716 13786 13728
rect 14366 13716 14372 13728
rect 13780 13688 14372 13716
rect 13780 13676 13786 13688
rect 14366 13676 14372 13688
rect 14424 13716 14430 13728
rect 14918 13716 14924 13728
rect 14424 13688 14924 13716
rect 14424 13676 14430 13688
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 1489 13515 1547 13521
rect 1489 13512 1501 13515
rect 860 13484 1501 13512
rect 860 13385 888 13484
rect 1489 13481 1501 13484
rect 1535 13512 1547 13515
rect 2498 13512 2504 13524
rect 1535 13484 2504 13512
rect 1535 13481 1547 13484
rect 1489 13475 1547 13481
rect 2498 13472 2504 13484
rect 2556 13472 2562 13524
rect 2869 13515 2927 13521
rect 2869 13481 2881 13515
rect 2915 13512 2927 13515
rect 2958 13512 2964 13524
rect 2915 13484 2964 13512
rect 2915 13481 2927 13484
rect 2869 13475 2927 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 4430 13472 4436 13524
rect 4488 13472 4494 13524
rect 8588 13484 12434 13512
rect 1121 13447 1179 13453
rect 1121 13413 1133 13447
rect 1167 13413 1179 13447
rect 1949 13447 2007 13453
rect 1949 13444 1961 13447
rect 1121 13407 1179 13413
rect 1412 13416 1961 13444
rect 845 13379 903 13385
rect 845 13345 857 13379
rect 891 13345 903 13379
rect 845 13339 903 13345
rect 1029 13379 1087 13385
rect 1029 13345 1041 13379
rect 1075 13376 1087 13379
rect 1136 13376 1164 13407
rect 1412 13385 1440 13416
rect 1949 13413 1961 13416
rect 1995 13413 2007 13447
rect 1949 13407 2007 13413
rect 8588 13388 8616 13484
rect 8938 13404 8944 13456
rect 8996 13444 9002 13456
rect 10321 13447 10379 13453
rect 8996 13416 9812 13444
rect 8996 13404 9002 13416
rect 1075 13348 1164 13376
rect 1397 13379 1455 13385
rect 1075 13345 1087 13348
rect 1029 13339 1087 13345
rect 1397 13345 1409 13379
rect 1443 13345 1455 13379
rect 1397 13339 1455 13345
rect 1670 13336 1676 13388
rect 1728 13336 1734 13388
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 5994 13336 6000 13388
rect 6052 13376 6058 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6052 13348 6745 13376
rect 6052 13336 6058 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 6917 13379 6975 13385
rect 6917 13345 6929 13379
rect 6963 13376 6975 13379
rect 7282 13376 7288 13388
rect 6963 13348 7288 13376
rect 6963 13345 6975 13348
rect 6917 13339 6975 13345
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 8478 13336 8484 13388
rect 8536 13336 8542 13388
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 9784 13385 9812 13416
rect 10321 13413 10333 13447
rect 10367 13444 10379 13447
rect 11210 13447 11268 13453
rect 11210 13444 11222 13447
rect 10367 13416 11222 13444
rect 10367 13413 10379 13416
rect 10321 13407 10379 13413
rect 11210 13413 11222 13416
rect 11256 13413 11268 13447
rect 11210 13407 11268 13413
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9769 13379 9827 13385
rect 9079 13348 9720 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 1121 13311 1179 13317
rect 1121 13277 1133 13311
rect 1167 13277 1179 13311
rect 1121 13271 1179 13277
rect 1305 13311 1363 13317
rect 1305 13277 1317 13311
rect 1351 13308 1363 13311
rect 1688 13308 1716 13336
rect 1351 13280 1716 13308
rect 1351 13277 1363 13280
rect 1305 13271 1363 13277
rect 1136 13240 1164 13271
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 1912 13280 2513 13308
rect 1912 13268 1918 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 3326 13308 3332 13320
rect 2648 13280 3332 13308
rect 2648 13268 2654 13280
rect 3326 13268 3332 13280
rect 3384 13308 3390 13320
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3384 13280 3433 13308
rect 3384 13268 3390 13280
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 8202 13308 8208 13320
rect 8159 13280 8208 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 8496 13308 8524 13336
rect 9122 13308 9128 13320
rect 8496 13280 9128 13308
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 9692 13308 9720 13348
rect 9769 13345 9781 13379
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10502 13336 10508 13388
rect 10560 13336 10566 13388
rect 10781 13379 10839 13385
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 11606 13376 11612 13388
rect 10827 13348 11612 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 10686 13308 10692 13320
rect 9692 13280 10692 13308
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 12406 13308 12434 13484
rect 15102 13472 15108 13524
rect 15160 13512 15166 13524
rect 15160 13484 17632 13512
rect 15160 13472 15166 13484
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 12618 13444 12624 13456
rect 12575 13416 12624 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 12710 13404 12716 13456
rect 12768 13453 12774 13456
rect 12768 13447 12787 13453
rect 12775 13413 12787 13447
rect 15194 13444 15200 13456
rect 12768 13407 12787 13413
rect 12912 13416 15200 13444
rect 12768 13404 12774 13407
rect 12912 13308 12940 13416
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 15749 13447 15807 13453
rect 15749 13413 15761 13447
rect 15795 13444 15807 13447
rect 15795 13416 17540 13444
rect 15795 13413 15807 13416
rect 15749 13407 15807 13413
rect 17512 13388 17540 13416
rect 13906 13336 13912 13388
rect 13964 13336 13970 13388
rect 13998 13336 14004 13388
rect 14056 13376 14062 13388
rect 14165 13379 14223 13385
rect 14165 13376 14177 13379
rect 14056 13348 14177 13376
rect 14056 13336 14062 13348
rect 14165 13345 14177 13348
rect 14211 13345 14223 13379
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 14165 13339 14223 13345
rect 15304 13348 15485 13376
rect 12406 13280 12940 13308
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13308 13323 13311
rect 13538 13308 13544 13320
rect 13311 13280 13544 13308
rect 13311 13277 13323 13280
rect 13265 13271 13323 13277
rect 2314 13240 2320 13252
rect 1136 13212 2320 13240
rect 2314 13200 2320 13212
rect 2372 13200 2378 13252
rect 10778 13240 10784 13252
rect 9968 13212 10784 13240
rect 1026 13132 1032 13184
rect 1084 13132 1090 13184
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13172 6883 13175
rect 6914 13172 6920 13184
rect 6871 13144 6920 13172
rect 6871 13141 6883 13144
rect 6825 13135 6883 13141
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 8757 13175 8815 13181
rect 8757 13172 8769 13175
rect 8720 13144 8769 13172
rect 8720 13132 8726 13144
rect 8757 13141 8769 13144
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 8846 13132 8852 13184
rect 8904 13132 8910 13184
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9968 13181 9996 13212
rect 10778 13200 10784 13212
rect 10836 13200 10842 13252
rect 12897 13243 12955 13249
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 13004 13240 13032 13271
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 15304 13249 15332 13348
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 16942 13336 16948 13388
rect 17000 13336 17006 13388
rect 17494 13336 17500 13388
rect 17552 13336 17558 13388
rect 17604 13376 17632 13484
rect 18138 13472 18144 13524
rect 18196 13472 18202 13524
rect 18509 13379 18567 13385
rect 18509 13376 18521 13379
rect 17604 13348 18521 13376
rect 18509 13345 18521 13348
rect 18555 13345 18567 13379
rect 18509 13339 18567 13345
rect 18598 13268 18604 13320
rect 18656 13268 18662 13320
rect 12943 13212 13032 13240
rect 15289 13243 15347 13249
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 15289 13209 15301 13243
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9732 13144 9965 13172
rect 9732 13132 9738 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 10689 13175 10747 13181
rect 10689 13141 10701 13175
rect 10735 13172 10747 13175
rect 11146 13172 11152 13184
rect 10735 13144 11152 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12345 13175 12403 13181
rect 12345 13172 12357 13175
rect 12124 13144 12357 13172
rect 12124 13132 12130 13144
rect 12345 13141 12357 13144
rect 12391 13141 12403 13175
rect 12345 13135 12403 13141
rect 12526 13132 12532 13184
rect 12584 13172 12590 13184
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 12584 13144 12725 13172
rect 12584 13132 12590 13144
rect 12713 13141 12725 13144
rect 12759 13172 12771 13175
rect 13722 13172 13728 13184
rect 12759 13144 13728 13172
rect 12759 13141 12771 13144
rect 12713 13135 12771 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 16114 13132 16120 13184
rect 16172 13132 16178 13184
rect 18782 13132 18788 13184
rect 18840 13132 18846 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 1854 12928 1860 12980
rect 1912 12968 1918 12980
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 1912 12940 3249 12968
rect 1912 12928 1918 12940
rect 3237 12937 3249 12940
rect 3283 12937 3295 12971
rect 3237 12931 3295 12937
rect 8021 12971 8079 12977
rect 8021 12937 8033 12971
rect 8067 12937 8079 12971
rect 8021 12931 8079 12937
rect 3697 12903 3755 12909
rect 3697 12869 3709 12903
rect 3743 12900 3755 12903
rect 7190 12900 7196 12912
rect 3743 12872 7196 12900
rect 3743 12869 3755 12872
rect 3697 12863 3755 12869
rect 7190 12860 7196 12872
rect 7248 12860 7254 12912
rect 8036 12900 8064 12931
rect 8202 12928 8208 12980
rect 8260 12928 8266 12980
rect 8754 12968 8760 12980
rect 8312 12940 8760 12968
rect 8312 12900 8340 12940
rect 8754 12928 8760 12940
rect 8812 12968 8818 12980
rect 9214 12968 9220 12980
rect 8812 12940 9220 12968
rect 8812 12928 8818 12940
rect 9214 12928 9220 12940
rect 9272 12968 9278 12980
rect 9272 12940 9536 12968
rect 9272 12928 9278 12940
rect 8036 12872 8340 12900
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 1026 12792 1032 12844
rect 1084 12792 1090 12844
rect 3326 12792 3332 12844
rect 3384 12792 3390 12844
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12832 7987 12835
rect 8496 12832 8524 12860
rect 7975 12804 8524 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3108 12736 3464 12764
rect 3108 12724 3114 12736
rect 2808 12699 2866 12705
rect 2808 12665 2820 12699
rect 2854 12696 2866 12699
rect 3142 12696 3148 12708
rect 2854 12668 3148 12696
rect 2854 12665 2866 12668
rect 2808 12659 2866 12665
rect 3142 12656 3148 12668
rect 3200 12656 3206 12708
rect 3234 12656 3240 12708
rect 3292 12656 3298 12708
rect 3436 12696 3464 12736
rect 3510 12724 3516 12776
rect 3568 12724 3574 12776
rect 7098 12724 7104 12776
rect 7156 12724 7162 12776
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7650 12764 7656 12776
rect 7340 12736 7656 12764
rect 7340 12724 7346 12736
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 8478 12724 8484 12776
rect 8536 12724 8542 12776
rect 9508 12764 9536 12940
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10560 12940 10977 12968
rect 10560 12928 10566 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11072 12940 13032 12968
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 11072 12900 11100 12940
rect 12066 12900 12072 12912
rect 10744 12872 11100 12900
rect 11716 12872 12072 12900
rect 10744 12860 10750 12872
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11388 12804 11652 12832
rect 11388 12792 11394 12804
rect 11624 12776 11652 12804
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 9508 12736 10977 12764
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11241 12767 11299 12773
rect 11241 12764 11253 12767
rect 11204 12736 11253 12764
rect 11204 12724 11210 12736
rect 11241 12733 11253 12736
rect 11287 12764 11299 12767
rect 11514 12764 11520 12776
rect 11287 12736 11520 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 3970 12696 3976 12708
rect 3436 12668 3976 12696
rect 3970 12656 3976 12668
rect 4028 12696 4034 12708
rect 6454 12696 6460 12708
rect 4028 12668 6460 12696
rect 4028 12656 4034 12668
rect 1578 12588 1584 12640
rect 1636 12588 1642 12640
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12628 1731 12631
rect 2590 12628 2596 12640
rect 1719 12600 2596 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 5828 12637 5856 12668
rect 6454 12656 6460 12668
rect 6512 12696 6518 12708
rect 8496 12696 8524 12724
rect 6512 12668 8524 12696
rect 8748 12699 8806 12705
rect 6512 12656 6518 12668
rect 8748 12665 8760 12699
rect 8794 12696 8806 12699
rect 8846 12696 8852 12708
rect 8794 12668 8852 12696
rect 8794 12665 8806 12668
rect 8748 12659 8806 12665
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 11716 12696 11744 12872
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 12124 12872 12940 12900
rect 12124 12860 12130 12872
rect 12912 12844 12940 12872
rect 12268 12804 12848 12832
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 12069 12767 12127 12773
rect 12069 12764 12081 12767
rect 11839 12736 12081 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 12069 12733 12081 12736
rect 12115 12733 12127 12767
rect 12069 12727 12127 12733
rect 12158 12724 12164 12776
rect 12216 12764 12222 12776
rect 12268 12773 12296 12804
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12216 12736 12265 12764
rect 12216 12724 12222 12736
rect 12253 12733 12265 12736
rect 12299 12733 12311 12767
rect 12253 12727 12311 12733
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 11164 12668 11744 12696
rect 12360 12696 12388 12727
rect 12618 12724 12624 12776
rect 12676 12724 12682 12776
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 12820 12764 12848 12804
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13004 12832 13032 12940
rect 13078 12928 13084 12980
rect 13136 12928 13142 12980
rect 13998 12928 14004 12980
rect 14056 12928 14062 12980
rect 18414 12928 18420 12980
rect 18472 12968 18478 12980
rect 18598 12968 18604 12980
rect 18472 12940 18604 12968
rect 18472 12928 18478 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 13265 12903 13323 12909
rect 13265 12869 13277 12903
rect 13311 12900 13323 12903
rect 16666 12900 16672 12912
rect 13311 12872 16672 12900
rect 13311 12869 13323 12872
rect 13265 12863 13323 12869
rect 16666 12860 16672 12872
rect 16724 12860 16730 12912
rect 14182 12832 14188 12844
rect 13004 12804 14188 12832
rect 14182 12792 14188 12804
rect 14240 12792 14246 12844
rect 14458 12792 14464 12844
rect 14516 12792 14522 12844
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 14918 12832 14924 12844
rect 14783 12804 14924 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 15286 12792 15292 12844
rect 15344 12832 15350 12844
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 15344 12804 17049 12832
rect 15344 12792 15350 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12820 12736 13093 12764
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 13814 12724 13820 12776
rect 13872 12724 13878 12776
rect 13909 12767 13967 12773
rect 13909 12733 13921 12767
rect 13955 12733 13967 12767
rect 13909 12727 13967 12733
rect 12636 12696 12664 12724
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12360 12668 12817 12696
rect 5813 12631 5871 12637
rect 5813 12597 5825 12631
rect 5859 12597 5871 12631
rect 5813 12591 5871 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 11164 12637 11192 12668
rect 12805 12665 12817 12668
rect 12851 12665 12863 12699
rect 13633 12699 13691 12705
rect 13633 12696 13645 12699
rect 12805 12659 12863 12665
rect 12912 12668 13645 12696
rect 9861 12631 9919 12637
rect 9861 12628 9873 12631
rect 9732 12600 9873 12628
rect 9732 12588 9738 12600
rect 9861 12597 9873 12600
rect 9907 12597 9919 12631
rect 9861 12591 9919 12597
rect 11149 12631 11207 12637
rect 11149 12597 11161 12631
rect 11195 12597 11207 12631
rect 11149 12591 11207 12597
rect 11422 12588 11428 12640
rect 11480 12628 11486 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 11480 12600 11621 12628
rect 11480 12588 11486 12600
rect 11609 12597 11621 12600
rect 11655 12597 11667 12631
rect 11609 12591 11667 12597
rect 12434 12588 12440 12640
rect 12492 12588 12498 12640
rect 12526 12588 12532 12640
rect 12584 12628 12590 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12584 12600 12633 12628
rect 12584 12588 12590 12600
rect 12621 12597 12633 12600
rect 12667 12628 12679 12631
rect 12912 12628 12940 12668
rect 13633 12665 13645 12668
rect 13679 12665 13691 12699
rect 13924 12696 13952 12727
rect 14366 12724 14372 12776
rect 14424 12724 14430 12776
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 17304 12767 17362 12773
rect 16163 12736 16896 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 15102 12696 15108 12708
rect 13924 12668 15108 12696
rect 13633 12659 13691 12665
rect 15102 12656 15108 12668
rect 15160 12656 15166 12708
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 16540 12668 16773 12696
rect 16540 12656 16546 12668
rect 16761 12665 16773 12668
rect 16807 12665 16819 12699
rect 16761 12659 16819 12665
rect 16868 12640 16896 12736
rect 17304 12733 17316 12767
rect 17350 12764 17362 12767
rect 18782 12764 18788 12776
rect 17350 12736 18788 12764
rect 17350 12733 17362 12736
rect 17304 12727 17362 12733
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 12667 12600 12940 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 16850 12588 16856 12640
rect 16908 12628 16914 12640
rect 17494 12628 17500 12640
rect 16908 12600 17500 12628
rect 16908 12588 16914 12600
rect 17494 12588 17500 12600
rect 17552 12588 17558 12640
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 845 12427 903 12433
rect 845 12393 857 12427
rect 891 12424 903 12427
rect 1854 12424 1860 12436
rect 891 12396 1860 12424
rect 891 12393 903 12396
rect 845 12387 903 12393
rect 1854 12384 1860 12396
rect 1912 12424 1918 12436
rect 1912 12396 2452 12424
rect 1912 12384 1918 12396
rect 1578 12316 1584 12368
rect 1636 12356 1642 12368
rect 2424 12365 2452 12396
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4909 12427 4967 12433
rect 4909 12424 4921 12427
rect 4120 12396 4921 12424
rect 4120 12384 4126 12396
rect 4909 12393 4921 12396
rect 4955 12393 4967 12427
rect 4909 12387 4967 12393
rect 6822 12384 6828 12436
rect 6880 12384 6886 12436
rect 7944 12396 9076 12424
rect 1958 12359 2016 12365
rect 1958 12356 1970 12359
rect 1636 12328 1970 12356
rect 1636 12316 1642 12328
rect 1958 12325 1970 12328
rect 2004 12325 2016 12359
rect 1958 12319 2016 12325
rect 2409 12359 2467 12365
rect 2409 12325 2421 12359
rect 2455 12325 2467 12359
rect 2609 12359 2667 12365
rect 2609 12356 2621 12359
rect 2409 12319 2467 12325
rect 2516 12328 2621 12356
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 2516 12288 2544 12328
rect 2609 12325 2621 12328
rect 2655 12325 2667 12359
rect 2609 12319 2667 12325
rect 3988 12328 4660 12356
rect 3988 12297 4016 12328
rect 1728 12260 2544 12288
rect 3973 12291 4031 12297
rect 1728 12248 1734 12260
rect 3973 12257 3985 12291
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 3050 12220 3056 12232
rect 2280 12192 3056 12220
rect 2280 12180 2286 12192
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4172 12220 4200 12251
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 4632 12288 4660 12328
rect 4706 12316 4712 12368
rect 4764 12316 4770 12368
rect 5994 12356 6000 12368
rect 5368 12328 6000 12356
rect 4982 12288 4988 12300
rect 4632 12260 4988 12288
rect 4982 12248 4988 12260
rect 5040 12288 5046 12300
rect 5368 12297 5396 12328
rect 5994 12316 6000 12328
rect 6052 12316 6058 12368
rect 6914 12316 6920 12368
rect 6972 12316 6978 12368
rect 7374 12316 7380 12368
rect 7432 12316 7438 12368
rect 5353 12291 5411 12297
rect 5353 12288 5365 12291
rect 5040 12260 5365 12288
rect 5040 12248 5046 12260
rect 5353 12257 5365 12260
rect 5399 12257 5411 12291
rect 5534 12288 5540 12300
rect 5353 12251 5411 12257
rect 5460 12260 5540 12288
rect 5460 12220 5488 12260
rect 5534 12248 5540 12260
rect 5592 12288 5598 12300
rect 5810 12288 5816 12300
rect 5592 12260 5816 12288
rect 5592 12248 5598 12260
rect 5810 12248 5816 12260
rect 5868 12288 5874 12300
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 5868 12260 6469 12288
rect 5868 12248 5874 12260
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7193 12291 7251 12297
rect 7193 12288 7205 12291
rect 7156 12260 7205 12288
rect 7156 12248 7162 12260
rect 7193 12257 7205 12260
rect 7239 12257 7251 12291
rect 7193 12251 7251 12257
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 4172 12192 5488 12220
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7944 12220 7972 12396
rect 8478 12316 8484 12368
rect 8536 12356 8542 12368
rect 9048 12356 9076 12396
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 9548 12396 9597 12424
rect 9548 12384 9554 12396
rect 9585 12393 9597 12396
rect 9631 12393 9643 12427
rect 9585 12387 9643 12393
rect 8536 12328 8984 12356
rect 8536 12316 8542 12328
rect 8662 12248 8668 12300
rect 8720 12297 8726 12300
rect 8956 12297 8984 12328
rect 9048 12328 9628 12356
rect 9048 12297 9076 12328
rect 8720 12288 8732 12297
rect 8941 12291 8999 12297
rect 8720 12260 8765 12288
rect 8720 12251 8732 12260
rect 8941 12257 8953 12291
rect 8987 12257 8999 12291
rect 8941 12251 8999 12257
rect 9033 12291 9091 12297
rect 9033 12257 9045 12291
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 8720 12248 8726 12251
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 9180 12260 9321 12288
rect 9180 12248 9186 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9600 12288 9628 12328
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 11238 12356 11244 12368
rect 9732 12328 11244 12356
rect 9732 12316 9738 12328
rect 11238 12316 11244 12328
rect 11296 12356 11302 12368
rect 12345 12359 12403 12365
rect 12345 12356 12357 12359
rect 11296 12328 12357 12356
rect 11296 12316 11302 12328
rect 12345 12325 12357 12328
rect 12391 12325 12403 12359
rect 12345 12319 12403 12325
rect 13906 12316 13912 12368
rect 13964 12316 13970 12368
rect 9766 12288 9772 12300
rect 9600 12260 9772 12288
rect 9309 12251 9367 12257
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 11054 12248 11060 12300
rect 11112 12248 11118 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 6595 12192 7972 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 5169 12155 5227 12161
rect 5169 12152 5181 12155
rect 4908 12124 5181 12152
rect 2590 12044 2596 12096
rect 2648 12044 2654 12096
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 3142 12084 3148 12096
rect 2823 12056 3148 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12084 4491 12087
rect 4522 12084 4528 12096
rect 4479 12056 4528 12084
rect 4479 12053 4491 12056
rect 4433 12047 4491 12053
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 4908 12093 4936 12124
rect 5169 12121 5181 12124
rect 5215 12121 5227 12155
rect 11164 12152 11192 12251
rect 11422 12248 11428 12300
rect 11480 12248 11486 12300
rect 11514 12248 11520 12300
rect 11572 12288 11578 12300
rect 13630 12288 13636 12300
rect 11572 12260 13636 12288
rect 11572 12248 11578 12260
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 17310 12248 17316 12300
rect 17368 12248 17374 12300
rect 17494 12248 17500 12300
rect 17552 12248 17558 12300
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12220 11299 12223
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11287 12192 11621 12220
rect 11287 12189 11299 12192
rect 11241 12183 11299 12189
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12161 12223 12219 12229
rect 12161 12220 12173 12223
rect 12124 12192 12173 12220
rect 12124 12180 12130 12192
rect 12161 12189 12173 12192
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12526 12152 12532 12164
rect 11164 12124 12532 12152
rect 5169 12115 5227 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 4893 12087 4951 12093
rect 4893 12053 4905 12087
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 5077 12087 5135 12093
rect 5077 12053 5089 12087
rect 5123 12084 5135 12087
rect 5810 12084 5816 12096
rect 5123 12056 5816 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7340 12056 7573 12084
rect 7340 12044 7346 12056
rect 7561 12053 7573 12056
rect 7607 12084 7619 12087
rect 7650 12084 7656 12096
rect 7607 12056 7656 12084
rect 7607 12053 7619 12056
rect 7561 12047 7619 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 9214 12044 9220 12096
rect 9272 12044 9278 12096
rect 11422 12044 11428 12096
rect 11480 12044 11486 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 16485 12087 16543 12093
rect 16485 12084 16497 12087
rect 15068 12056 16497 12084
rect 15068 12044 15074 12056
rect 16485 12053 16497 12056
rect 16531 12053 16543 12087
rect 16485 12047 16543 12053
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 3142 11880 3148 11892
rect 2915 11852 3148 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3142 11840 3148 11852
rect 3200 11880 3206 11892
rect 3418 11880 3424 11892
rect 3200 11852 3424 11880
rect 3200 11840 3206 11852
rect 3418 11840 3424 11852
rect 3476 11880 3482 11892
rect 4062 11880 4068 11892
rect 3476 11852 4068 11880
rect 3476 11840 3482 11852
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4304 11852 4537 11880
rect 4304 11840 4310 11852
rect 4525 11849 4537 11852
rect 4571 11849 4583 11883
rect 4525 11843 4583 11849
rect 5077 11883 5135 11889
rect 5077 11849 5089 11883
rect 5123 11880 5135 11883
rect 5534 11880 5540 11892
rect 5123 11852 5540 11880
rect 5123 11849 5135 11852
rect 5077 11843 5135 11849
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 7006 11840 7012 11892
rect 7064 11840 7070 11892
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9674 11880 9680 11892
rect 9539 11852 9680 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 12345 11883 12403 11889
rect 12345 11849 12357 11883
rect 12391 11880 12403 11883
rect 12526 11880 12532 11892
rect 12391 11852 12532 11880
rect 12391 11849 12403 11852
rect 12345 11843 12403 11849
rect 12526 11840 12532 11852
rect 12584 11880 12590 11892
rect 12584 11852 12940 11880
rect 12584 11840 12590 11852
rect 2314 11772 2320 11824
rect 2372 11812 2378 11824
rect 2372 11784 3924 11812
rect 2372 11772 2378 11784
rect 2700 11753 2728 11784
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3234 11704 3240 11756
rect 3292 11704 3298 11756
rect 3896 11744 3924 11784
rect 3970 11772 3976 11824
rect 4028 11772 4034 11824
rect 4617 11815 4675 11821
rect 4617 11781 4629 11815
rect 4663 11812 4675 11815
rect 4706 11812 4712 11824
rect 4663 11784 4712 11812
rect 4663 11781 4675 11784
rect 4617 11775 4675 11781
rect 4632 11744 4660 11775
rect 4706 11772 4712 11784
rect 4764 11772 4770 11824
rect 3896 11716 4660 11744
rect 4982 11704 4988 11756
rect 5040 11704 5046 11756
rect 6454 11704 6460 11756
rect 6512 11704 6518 11756
rect 12802 11744 12808 11756
rect 12544 11716 12808 11744
rect 2961 11679 3019 11685
rect 2961 11645 2973 11679
rect 3007 11676 3019 11679
rect 3881 11679 3939 11685
rect 3881 11676 3893 11679
rect 3007 11648 3893 11676
rect 3007 11645 3019 11648
rect 2961 11639 3019 11645
rect 3881 11645 3893 11648
rect 3927 11676 3939 11679
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 3927 11648 4169 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11645 4307 11679
rect 5000 11676 5028 11704
rect 6641 11679 6699 11685
rect 5000 11648 6316 11676
rect 4249 11639 4307 11645
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11608 2743 11611
rect 3973 11611 4031 11617
rect 3973 11608 3985 11611
rect 2731 11580 3985 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 3973 11577 3985 11580
rect 4019 11577 4031 11611
rect 3973 11571 4031 11577
rect 4062 11568 4068 11620
rect 4120 11608 4126 11620
rect 4264 11608 4292 11639
rect 4120 11580 4292 11608
rect 4120 11568 4126 11580
rect 5994 11568 6000 11620
rect 6052 11608 6058 11620
rect 6190 11611 6248 11617
rect 6190 11608 6202 11611
rect 6052 11580 6202 11608
rect 6052 11568 6058 11580
rect 6190 11577 6202 11580
rect 6236 11577 6248 11611
rect 6288 11608 6316 11648
rect 6641 11645 6653 11679
rect 6687 11676 6699 11679
rect 7282 11676 7288 11688
rect 6687 11648 7288 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 10778 11636 10784 11688
rect 10836 11636 10842 11688
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 10962 11676 10968 11688
rect 10919 11648 10968 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11140 11679 11198 11685
rect 11140 11645 11152 11679
rect 11186 11676 11198 11679
rect 11422 11676 11428 11688
rect 11186 11648 11428 11676
rect 11186 11645 11198 11648
rect 11140 11639 11198 11645
rect 11422 11636 11428 11648
rect 11480 11636 11486 11688
rect 12544 11685 12572 11716
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 12529 11679 12587 11685
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 12710 11636 12716 11688
rect 12768 11636 12774 11688
rect 12912 11685 12940 11852
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 13872 11852 14289 11880
rect 13872 11840 13878 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 15197 11883 15255 11889
rect 15197 11849 15209 11883
rect 15243 11880 15255 11883
rect 15930 11880 15936 11892
rect 15243 11852 15936 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15930 11840 15936 11852
rect 15988 11840 15994 11892
rect 13262 11772 13268 11824
rect 13320 11812 13326 11824
rect 13320 11784 14596 11812
rect 13320 11772 13326 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11744 13231 11747
rect 13446 11744 13452 11756
rect 13219 11716 13452 11744
rect 13219 11713 13231 11716
rect 13173 11707 13231 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 13556 11716 14473 11744
rect 13556 11685 13584 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14568 11744 14596 11784
rect 16390 11744 16396 11756
rect 14568 11716 16396 11744
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13541 11679 13599 11685
rect 13541 11676 13553 11679
rect 13127 11648 13553 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13541 11645 13553 11648
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 6825 11611 6883 11617
rect 6825 11608 6837 11611
rect 6288 11580 6837 11608
rect 6190 11571 6248 11577
rect 6825 11577 6837 11580
rect 6871 11577 6883 11611
rect 12912 11608 12940 11639
rect 13630 11636 13636 11688
rect 13688 11676 13694 11688
rect 14568 11685 14596 11716
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 14001 11679 14059 11685
rect 14001 11676 14013 11679
rect 13688 11648 14013 11676
rect 13688 11636 13694 11648
rect 14001 11645 14013 11648
rect 14047 11645 14059 11679
rect 14369 11679 14427 11685
rect 14369 11676 14381 11679
rect 14001 11639 14059 11645
rect 14108 11648 14381 11676
rect 14108 11617 14136 11648
rect 14369 11645 14381 11648
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 13725 11611 13783 11617
rect 13725 11608 13737 11611
rect 12912 11580 13737 11608
rect 6825 11571 6883 11577
rect 13725 11577 13737 11580
rect 13771 11577 13783 11611
rect 14093 11611 14151 11617
rect 14093 11608 14105 11611
rect 13725 11571 13783 11577
rect 13832 11580 14105 11608
rect 10594 11500 10600 11552
rect 10652 11540 10658 11552
rect 12066 11540 12072 11552
rect 10652 11512 12072 11540
rect 10652 11500 10658 11512
rect 12066 11500 12072 11512
rect 12124 11540 12130 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 12124 11512 12265 11540
rect 12124 11500 12130 11512
rect 12253 11509 12265 11512
rect 12299 11509 12311 11543
rect 12253 11503 12311 11509
rect 12986 11500 12992 11552
rect 13044 11540 13050 11552
rect 13832 11540 13860 11580
rect 14093 11577 14105 11580
rect 14139 11577 14151 11611
rect 14093 11571 14151 11577
rect 14277 11611 14335 11617
rect 14277 11577 14289 11611
rect 14323 11608 14335 11611
rect 14568 11608 14596 11639
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14976 11648 15025 11676
rect 14976 11636 14982 11648
rect 15013 11645 15025 11648
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 15105 11679 15163 11685
rect 15105 11645 15117 11679
rect 15151 11645 15163 11679
rect 15105 11639 15163 11645
rect 15120 11608 15148 11639
rect 15194 11636 15200 11688
rect 15252 11676 15258 11688
rect 16301 11679 16359 11685
rect 16301 11676 16313 11679
rect 15252 11648 16313 11676
rect 15252 11636 15258 11648
rect 16301 11645 16313 11648
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16758 11636 16764 11688
rect 16816 11636 16822 11688
rect 14323 11580 14596 11608
rect 15028 11580 15148 11608
rect 14323 11577 14335 11580
rect 14277 11571 14335 11577
rect 15028 11552 15056 11580
rect 13044 11512 13860 11540
rect 13909 11543 13967 11549
rect 13044 11500 13050 11512
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14182 11540 14188 11552
rect 13955 11512 14188 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 15010 11500 15016 11552
rect 15068 11500 15074 11552
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 15381 11543 15439 11549
rect 15381 11540 15393 11543
rect 15344 11512 15393 11540
rect 15344 11500 15350 11512
rect 15381 11509 15393 11512
rect 15427 11509 15439 11543
rect 15381 11503 15439 11509
rect 15930 11500 15936 11552
rect 15988 11540 15994 11552
rect 16482 11540 16488 11552
rect 15988 11512 16488 11540
rect 15988 11500 15994 11512
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 2222 11336 2228 11348
rect 2056 11308 2228 11336
rect 2056 11268 2084 11308
rect 2222 11296 2228 11308
rect 2280 11296 2286 11348
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3421 11339 3479 11345
rect 3421 11336 3433 11339
rect 3292 11308 3433 11336
rect 3292 11296 3298 11308
rect 3421 11305 3433 11308
rect 3467 11305 3479 11339
rect 3421 11299 3479 11305
rect 4982 11296 4988 11348
rect 5040 11336 5046 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 5040 11308 5641 11336
rect 5040 11296 5046 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5629 11299 5687 11305
rect 5994 11296 6000 11348
rect 6052 11296 6058 11348
rect 2056 11240 4292 11268
rect 2056 11209 2084 11240
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11169 2099 11203
rect 2041 11163 2099 11169
rect 2308 11203 2366 11209
rect 2308 11169 2320 11203
rect 2354 11200 2366 11203
rect 3970 11200 3976 11212
rect 2354 11172 3976 11200
rect 2354 11169 2366 11172
rect 2308 11163 2366 11169
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4264 11209 4292 11240
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 10410 11268 10416 11280
rect 8628 11240 8984 11268
rect 8628 11228 8634 11240
rect 4522 11209 4528 11212
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4516 11200 4528 11209
rect 4483 11172 4528 11200
rect 4249 11163 4307 11169
rect 4516 11163 4528 11172
rect 4522 11160 4528 11163
rect 4580 11160 4586 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 8956 11209 8984 11240
rect 9140 11240 10416 11268
rect 9140 11209 9168 11240
rect 9600 11212 9628 11240
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 13078 11228 13084 11280
rect 13136 11228 13142 11280
rect 17402 11268 17408 11280
rect 15120 11240 17408 11268
rect 15120 11212 15148 11240
rect 17402 11228 17408 11240
rect 17460 11268 17466 11280
rect 17460 11240 17724 11268
rect 17460 11228 17466 11240
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9125 11203 9183 11209
rect 9125 11169 9137 11203
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 8772 11132 8800 11163
rect 9140 11132 9168 11163
rect 9306 11160 9312 11212
rect 9364 11160 9370 11212
rect 9398 11160 9404 11212
rect 9456 11160 9462 11212
rect 9582 11160 9588 11212
rect 9640 11160 9646 11212
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 13262 11160 13268 11212
rect 13320 11160 13326 11212
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 15102 11200 15108 11212
rect 14875 11172 15108 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 17696 11209 17724 11240
rect 17862 11228 17868 11280
rect 17920 11268 17926 11280
rect 17920 11240 18078 11268
rect 17920 11228 17926 11240
rect 16577 11203 16635 11209
rect 16577 11200 16589 11203
rect 16448 11172 16589 11200
rect 16448 11160 16454 11172
rect 16577 11169 16589 11172
rect 16623 11200 16635 11203
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 16623 11172 17141 11200
rect 16623 11169 16635 11172
rect 16577 11163 16635 11169
rect 17129 11169 17141 11172
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 8772 11104 9168 11132
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11132 14151 11135
rect 14182 11132 14188 11144
rect 14139 11104 14188 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 14921 11095 14979 11101
rect 8849 11067 8907 11073
rect 8849 11033 8861 11067
rect 8895 11064 8907 11067
rect 8938 11064 8944 11076
rect 8895 11036 8944 11064
rect 8895 11033 8907 11036
rect 8849 11027 8907 11033
rect 8938 11024 8944 11036
rect 8996 11024 9002 11076
rect 9217 11067 9275 11073
rect 9217 11033 9229 11067
rect 9263 11064 9275 11067
rect 9306 11064 9312 11076
rect 9263 11036 9312 11064
rect 9263 11033 9275 11036
rect 9217 11027 9275 11033
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 9493 11067 9551 11073
rect 9493 11033 9505 11067
rect 9539 11064 9551 11067
rect 10226 11064 10232 11076
rect 9539 11036 10232 11064
rect 9539 11033 9551 11036
rect 9493 11027 9551 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 14936 11064 14964 11095
rect 16666 11092 16672 11144
rect 16724 11092 16730 11144
rect 17218 11064 17224 11076
rect 14936 11036 17224 11064
rect 17218 11024 17224 11036
rect 17276 11024 17282 11076
rect 16945 10999 17003 11005
rect 16945 10965 16957 10999
rect 16991 10996 17003 10999
rect 17402 10996 17408 11008
rect 16991 10968 17408 10996
rect 16991 10965 17003 10968
rect 16945 10959 17003 10965
rect 17402 10956 17408 10968
rect 17460 10956 17466 11008
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 13078 10752 13084 10804
rect 13136 10792 13142 10804
rect 14918 10792 14924 10804
rect 13136 10764 14924 10792
rect 13136 10752 13142 10764
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 10962 10724 10968 10736
rect 10827 10696 10968 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 16482 10724 16488 10736
rect 14108 10696 16488 10724
rect 10137 10659 10195 10665
rect 10137 10625 10149 10659
rect 10183 10656 10195 10659
rect 10183 10628 10824 10656
rect 10183 10625 10195 10628
rect 10137 10619 10195 10625
rect 10796 10600 10824 10628
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 14108 10600 14136 10696
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 14366 10656 14372 10668
rect 14292 10628 14372 10656
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 7984 10560 8401 10588
rect 7984 10548 7990 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 9582 10588 9588 10600
rect 8619 10560 9588 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 9582 10548 9588 10560
rect 9640 10588 9646 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9640 10560 10057 10588
rect 9640 10548 9646 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10594 10548 10600 10600
rect 10652 10548 10658 10600
rect 10778 10548 10784 10600
rect 10836 10548 10842 10600
rect 12710 10548 12716 10600
rect 12768 10588 12774 10600
rect 13262 10588 13268 10600
rect 12768 10560 13268 10588
rect 12768 10548 12774 10560
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 14090 10548 14096 10600
rect 14148 10548 14154 10600
rect 14292 10597 14320 10628
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 15010 10656 15016 10668
rect 14424 10628 15016 10656
rect 14424 10616 14430 10628
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 14277 10591 14335 10597
rect 14277 10557 14289 10591
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14829 10591 14887 10597
rect 14829 10557 14841 10591
rect 14875 10588 14887 10591
rect 15194 10588 15200 10600
rect 14875 10560 15200 10588
rect 14875 10557 14887 10560
rect 14829 10551 14887 10557
rect 13280 10492 13952 10520
rect 13280 10464 13308 10492
rect 8481 10455 8539 10461
rect 8481 10421 8493 10455
rect 8527 10452 8539 10455
rect 9674 10452 9680 10464
rect 8527 10424 9680 10452
rect 8527 10421 8539 10424
rect 8481 10415 8539 10421
rect 9674 10412 9680 10424
rect 9732 10412 9738 10464
rect 13262 10412 13268 10464
rect 13320 10412 13326 10464
rect 13354 10412 13360 10464
rect 13412 10412 13418 10464
rect 13924 10452 13952 10492
rect 13998 10480 14004 10532
rect 14056 10520 14062 10532
rect 14369 10523 14427 10529
rect 14369 10520 14381 10523
rect 14056 10492 14381 10520
rect 14056 10480 14062 10492
rect 14369 10489 14381 10492
rect 14415 10489 14427 10523
rect 14568 10520 14596 10551
rect 15194 10548 15200 10560
rect 15252 10548 15258 10600
rect 16390 10548 16396 10600
rect 16448 10548 16454 10600
rect 16574 10548 16580 10600
rect 16632 10548 16638 10600
rect 17037 10591 17095 10597
rect 17037 10557 17049 10591
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 14921 10523 14979 10529
rect 14921 10520 14933 10523
rect 14568 10492 14933 10520
rect 14369 10483 14427 10489
rect 14921 10489 14933 10492
rect 14967 10520 14979 10523
rect 15102 10520 15108 10532
rect 14967 10492 15108 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 16408 10520 16436 10548
rect 17052 10520 17080 10551
rect 17218 10548 17224 10600
rect 17276 10548 17282 10600
rect 16408 10492 17080 10520
rect 18046 10480 18052 10532
rect 18104 10480 18110 10532
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13924 10424 14197 10452
rect 14185 10421 14197 10424
rect 14231 10452 14243 10455
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 14231 10424 14749 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 14737 10415 14795 10421
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11204 10220 11376 10248
rect 11204 10208 11210 10220
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 9640 10152 9720 10180
rect 9640 10140 9646 10152
rect 9692 10121 9720 10152
rect 9858 10140 9864 10192
rect 9916 10140 9922 10192
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 10836 10152 11284 10180
rect 10836 10140 10842 10152
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10275 10115 10333 10121
rect 10275 10112 10287 10115
rect 9723 10084 10287 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10275 10081 10287 10084
rect 10321 10081 10333 10115
rect 10275 10075 10333 10081
rect 10410 10072 10416 10124
rect 10468 10072 10474 10124
rect 10502 10072 10508 10124
rect 10560 10072 10566 10124
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 10870 10112 10876 10124
rect 10643 10084 10876 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 10962 10072 10968 10124
rect 11020 10072 11026 10124
rect 11256 10121 11284 10152
rect 11348 10121 11376 10220
rect 13446 10208 13452 10260
rect 13504 10248 13510 10260
rect 16669 10251 16727 10257
rect 13504 10220 14780 10248
rect 13504 10208 13510 10220
rect 13354 10140 13360 10192
rect 13412 10180 13418 10192
rect 13412 10152 14320 10180
rect 13412 10140 13418 10152
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10081 11207 10115
rect 11149 10075 11207 10081
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 11333 10115 11391 10121
rect 11333 10081 11345 10115
rect 11379 10081 11391 10115
rect 11333 10075 11391 10081
rect 13817 10115 13875 10121
rect 13817 10081 13829 10115
rect 13863 10081 13875 10115
rect 13817 10075 13875 10081
rect 14001 10115 14059 10121
rect 14001 10081 14013 10115
rect 14047 10112 14059 10115
rect 14090 10112 14096 10124
rect 14047 10084 14096 10112
rect 14047 10081 14059 10084
rect 14001 10075 14059 10081
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 10686 10044 10692 10056
rect 10183 10016 10692 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 10042 9936 10048 9988
rect 10100 9936 10106 9988
rect 10980 9976 11008 10072
rect 11164 10044 11192 10075
rect 11164 10016 11376 10044
rect 11348 9988 11376 10016
rect 10244 9948 11008 9976
rect 10134 9868 10140 9920
rect 10192 9908 10198 9920
rect 10244 9908 10272 9948
rect 11330 9936 11336 9988
rect 11388 9936 11394 9988
rect 12986 9936 12992 9988
rect 13044 9976 13050 9988
rect 13832 9976 13860 10075
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 14292 10121 14320 10152
rect 14752 10121 14780 10220
rect 16669 10217 16681 10251
rect 16715 10248 16727 10251
rect 18046 10248 18052 10260
rect 16715 10220 18052 10248
rect 16715 10217 16727 10220
rect 16669 10211 16727 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 15194 10140 15200 10192
rect 15252 10180 15258 10192
rect 16301 10183 16359 10189
rect 16301 10180 16313 10183
rect 15252 10152 16313 10180
rect 15252 10140 15258 10152
rect 16301 10149 16313 10152
rect 16347 10149 16359 10183
rect 16301 10143 16359 10149
rect 14277 10115 14335 10121
rect 14277 10081 14289 10115
rect 14323 10081 14335 10115
rect 14277 10075 14335 10081
rect 14553 10115 14611 10121
rect 14553 10081 14565 10115
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 14737 10115 14795 10121
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 13964 10016 14473 10044
rect 13964 10004 13970 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14568 10044 14596 10075
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15013 10115 15071 10121
rect 15013 10112 15025 10115
rect 14976 10084 15025 10112
rect 14976 10072 14982 10084
rect 15013 10081 15025 10084
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 15286 10072 15292 10124
rect 15344 10072 15350 10124
rect 16114 10072 16120 10124
rect 16172 10112 16178 10124
rect 16485 10115 16543 10121
rect 16485 10112 16497 10115
rect 16172 10084 16497 10112
rect 16172 10072 16178 10084
rect 16485 10081 16497 10084
rect 16531 10081 16543 10115
rect 16485 10075 16543 10081
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10081 16819 10115
rect 16761 10075 16819 10081
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 14568 10016 14841 10044
rect 14461 10007 14519 10013
rect 14829 10013 14841 10016
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 16574 10004 16580 10056
rect 16632 10044 16638 10056
rect 16776 10044 16804 10075
rect 17402 10072 17408 10124
rect 17460 10072 17466 10124
rect 17862 10044 17868 10056
rect 16632 10016 17868 10044
rect 16632 10004 16638 10016
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 14369 9979 14427 9985
rect 13044 9948 14228 9976
rect 13044 9936 13050 9948
rect 10192 9880 10272 9908
rect 10192 9868 10198 9880
rect 10778 9868 10784 9920
rect 10836 9868 10842 9920
rect 11606 9868 11612 9920
rect 11664 9868 11670 9920
rect 13906 9868 13912 9920
rect 13964 9868 13970 9920
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 14200 9908 14228 9948
rect 14369 9945 14381 9979
rect 14415 9976 14427 9979
rect 15286 9976 15292 9988
rect 14415 9948 15292 9976
rect 14415 9945 14427 9948
rect 14369 9939 14427 9945
rect 15286 9936 15292 9948
rect 15344 9976 15350 9988
rect 17221 9979 17279 9985
rect 17221 9976 17233 9979
rect 15344 9948 17233 9976
rect 15344 9936 15350 9948
rect 17221 9945 17233 9948
rect 17267 9945 17279 9979
rect 17221 9939 17279 9945
rect 16114 9908 16120 9920
rect 14200 9880 16120 9908
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10686 9704 10692 9716
rect 9732 9676 10692 9704
rect 9732 9664 9738 9676
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 12989 9707 13047 9713
rect 12989 9673 13001 9707
rect 13035 9704 13047 9707
rect 13170 9704 13176 9716
rect 13035 9676 13176 9704
rect 13035 9673 13047 9676
rect 12989 9667 13047 9673
rect 13170 9664 13176 9676
rect 13228 9704 13234 9716
rect 15286 9704 15292 9716
rect 13228 9676 15292 9704
rect 13228 9664 13234 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 8846 9596 8852 9648
rect 8904 9596 8910 9648
rect 9490 9636 9496 9648
rect 8956 9608 9496 9636
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9500 8907 9503
rect 8956 9500 8984 9608
rect 9490 9596 9496 9608
rect 9548 9596 9554 9648
rect 9766 9636 9772 9648
rect 9600 9608 9772 9636
rect 9600 9568 9628 9608
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 9876 9608 10609 9636
rect 9048 9540 9628 9568
rect 9677 9571 9735 9577
rect 9048 9509 9076 9540
rect 9677 9537 9689 9571
rect 9723 9568 9735 9571
rect 9876 9568 9904 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 13541 9639 13599 9645
rect 13541 9636 13553 9639
rect 10597 9599 10655 9605
rect 11348 9608 13553 9636
rect 9723 9540 9904 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10318 9568 10324 9580
rect 10008 9540 10324 9568
rect 10008 9528 10014 9540
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 11348 9568 11376 9608
rect 13541 9605 13553 9608
rect 13587 9605 13599 9639
rect 13814 9636 13820 9648
rect 13541 9599 13599 9605
rect 13740 9608 13820 9636
rect 10459 9540 11376 9568
rect 11885 9571 11943 9577
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 11885 9537 11897 9571
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12526 9568 12532 9580
rect 12207 9540 12532 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 8895 9472 8984 9500
rect 9033 9503 9091 9509
rect 8895 9469 8907 9472
rect 8849 9463 8907 9469
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9140 9432 9168 9463
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 10778 9500 10784 9512
rect 9631 9472 10784 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11900 9500 11928 9531
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 12986 9568 12992 9580
rect 12851 9540 12992 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 12986 9528 12992 9540
rect 13044 9528 13050 9580
rect 13262 9568 13268 9580
rect 13096 9540 13268 9568
rect 10928 9472 11928 9500
rect 12069 9503 12127 9509
rect 10928 9460 10934 9472
rect 12069 9469 12081 9503
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 9140 9404 9812 9432
rect 9214 9324 9220 9376
rect 9272 9324 9278 9376
rect 9784 9373 9812 9404
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10229 9435 10287 9441
rect 10229 9432 10241 9435
rect 10100 9404 10241 9432
rect 10100 9392 10106 9404
rect 10229 9401 10241 9404
rect 10275 9432 10287 9435
rect 10594 9432 10600 9444
rect 10275 9404 10600 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 12084 9432 12112 9463
rect 12250 9460 12256 9512
rect 12308 9460 12314 9512
rect 12360 9509 12480 9510
rect 12345 9503 12480 9509
rect 12345 9469 12357 9503
rect 12391 9500 12480 9503
rect 12894 9500 12900 9512
rect 12391 9482 12900 9500
rect 12391 9469 12403 9482
rect 12452 9472 12900 9482
rect 12345 9463 12403 9469
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13096 9509 13124 9540
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13740 9577 13768 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14274 9636 14280 9648
rect 13924 9608 14280 9636
rect 13924 9577 13952 9608
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15838 9636 15844 9648
rect 15252 9608 15844 9636
rect 15252 9596 15258 9608
rect 15838 9596 15844 9608
rect 15896 9596 15902 9648
rect 16022 9596 16028 9648
rect 16080 9636 16086 9648
rect 16393 9639 16451 9645
rect 16393 9636 16405 9639
rect 16080 9608 16405 9636
rect 16080 9596 16086 9608
rect 16393 9605 16405 9608
rect 16439 9636 16451 9639
rect 16942 9636 16948 9648
rect 16439 9608 16948 9636
rect 16439 9605 16451 9608
rect 16393 9599 16451 9605
rect 16942 9596 16948 9608
rect 17000 9596 17006 9648
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9537 13783 9571
rect 13725 9531 13783 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14090 9568 14096 9580
rect 14047 9540 14096 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 14182 9528 14188 9580
rect 14240 9568 14246 9580
rect 15746 9568 15752 9580
rect 14240 9540 15752 9568
rect 14240 9528 14246 9540
rect 15746 9528 15752 9540
rect 15804 9568 15810 9580
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 15804 9540 16865 9568
rect 15804 9528 15810 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17678 9568 17684 9580
rect 17083 9540 17684 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17678 9528 17684 9540
rect 17736 9528 17742 9580
rect 13081 9503 13139 9509
rect 13081 9469 13093 9503
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13357 9503 13415 9509
rect 13357 9469 13369 9503
rect 13403 9500 13415 9503
rect 13630 9500 13636 9512
rect 13403 9472 13636 9500
rect 13403 9469 13415 9472
rect 13357 9463 13415 9469
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 14369 9503 14427 9509
rect 14369 9469 14381 9503
rect 14415 9500 14427 9503
rect 15010 9500 15016 9512
rect 14415 9472 15016 9500
rect 14415 9469 14427 9472
rect 14369 9463 14427 9469
rect 13722 9432 13728 9444
rect 12084 9404 13728 9432
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 9769 9367 9827 9373
rect 9769 9333 9781 9367
rect 9815 9333 9827 9367
rect 9769 9327 9827 9333
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10318 9364 10324 9376
rect 10192 9336 10324 9364
rect 10192 9324 10198 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10778 9364 10784 9376
rect 10560 9336 10784 9364
rect 10560 9324 10566 9336
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 12529 9367 12587 9373
rect 12529 9333 12541 9367
rect 12575 9364 12587 9367
rect 12618 9364 12624 9376
rect 12575 9336 12624 9364
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 13078 9324 13084 9376
rect 13136 9364 13142 9376
rect 13173 9367 13231 9373
rect 13173 9364 13185 9367
rect 13136 9336 13185 9364
rect 13136 9324 13142 9336
rect 13173 9333 13185 9336
rect 13219 9333 13231 9367
rect 13173 9327 13231 9333
rect 13630 9324 13636 9376
rect 13688 9364 13694 9376
rect 13833 9364 13861 9463
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15838 9460 15844 9512
rect 15896 9460 15902 9512
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16574 9500 16580 9512
rect 16071 9472 16580 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16574 9460 16580 9472
rect 16632 9460 16638 9512
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 14516 9404 14565 9432
rect 14516 9392 14522 9404
rect 14553 9401 14565 9404
rect 14599 9432 14611 9435
rect 15933 9435 15991 9441
rect 15933 9432 15945 9435
rect 14599 9404 15945 9432
rect 14599 9401 14611 9404
rect 14553 9395 14611 9401
rect 15933 9401 15945 9404
rect 15979 9401 15991 9435
rect 15933 9395 15991 9401
rect 13688 9336 13861 9364
rect 13688 9324 13694 9336
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 15010 9324 15016 9376
rect 15068 9364 15074 9376
rect 16114 9364 16120 9376
rect 15068 9336 16120 9364
rect 15068 9324 15074 9336
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16482 9324 16488 9376
rect 16540 9364 16546 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16540 9336 16773 9364
rect 16540 9324 16546 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10410 9160 10416 9172
rect 10183 9132 10416 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 11330 9160 11336 9172
rect 10520 9132 11336 9160
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 10520 9092 10548 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 12894 9120 12900 9172
rect 12952 9120 12958 9172
rect 13630 9120 13636 9172
rect 13688 9120 13694 9172
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 13780 9132 15485 9160
rect 13780 9120 13786 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 16022 9160 16028 9172
rect 15473 9123 15531 9129
rect 15672 9132 16028 9160
rect 9456 9064 10548 9092
rect 11057 9095 11115 9101
rect 9456 9052 9462 9064
rect 11057 9061 11069 9095
rect 11103 9092 11115 9095
rect 11238 9092 11244 9104
rect 11103 9064 11244 9092
rect 11103 9061 11115 9064
rect 11057 9055 11115 9061
rect 11238 9052 11244 9064
rect 11296 9052 11302 9104
rect 14458 9092 14464 9104
rect 13188 9064 14464 9092
rect 13188 9036 13216 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 9214 8984 9220 9036
rect 9272 8984 9278 9036
rect 10045 9027 10103 9033
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10318 9024 10324 9036
rect 10091 8996 10324 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 13078 8984 13084 9036
rect 13136 8984 13142 9036
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 9024 13875 9027
rect 14182 9024 14188 9036
rect 13863 8996 14188 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14424 8996 14565 9024
rect 14424 8984 14430 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 9508 8888 9536 8919
rect 13262 8916 13268 8968
rect 13320 8916 13326 8968
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 13538 8956 13544 8968
rect 13403 8928 13544 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 13909 8959 13967 8965
rect 13909 8956 13921 8959
rect 13780 8928 13921 8956
rect 13780 8916 13786 8928
rect 13909 8925 13921 8928
rect 13955 8925 13967 8959
rect 13909 8919 13967 8925
rect 13998 8916 14004 8968
rect 14056 8916 14062 8968
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 14458 8956 14464 8968
rect 14139 8928 14464 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 14660 8956 14688 8987
rect 14734 8984 14740 9036
rect 14792 8984 14798 9036
rect 14921 9027 14979 9033
rect 14921 8993 14933 9027
rect 14967 9024 14979 9027
rect 15378 9024 15384 9036
rect 14967 8996 15384 9024
rect 14967 8993 14979 8996
rect 14921 8987 14979 8993
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15672 9033 15700 9132
rect 16022 9120 16028 9132
rect 16080 9120 16086 9172
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 16574 9160 16580 9172
rect 16264 9132 16580 9160
rect 16264 9120 16270 9132
rect 16574 9120 16580 9132
rect 16632 9120 16638 9172
rect 17494 9120 17500 9172
rect 17552 9120 17558 9172
rect 17678 9120 17684 9172
rect 17736 9160 17742 9172
rect 18230 9160 18236 9172
rect 17736 9132 18236 9160
rect 17736 9120 17742 9132
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18046 9092 18052 9104
rect 17880 9064 18052 9092
rect 15657 9027 15715 9033
rect 15657 8993 15669 9027
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16022 9024 16028 9036
rect 15979 8996 16028 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 15286 8956 15292 8968
rect 14660 8928 15292 8956
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15856 8956 15884 8987
rect 16022 8984 16028 8996
rect 16080 8984 16086 9036
rect 16482 8984 16488 9036
rect 16540 8984 16546 9036
rect 16942 8984 16948 9036
rect 17000 8984 17006 9036
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17460 8996 17601 9024
rect 17460 8984 17466 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 17678 8984 17684 9036
rect 17736 8984 17742 9036
rect 17770 8984 17776 9036
rect 17828 9024 17834 9036
rect 17880 9033 17908 9064
rect 18046 9052 18052 9064
rect 18104 9052 18110 9104
rect 17865 9027 17923 9033
rect 17865 9024 17877 9027
rect 17828 8996 17877 9024
rect 17828 8984 17834 8996
rect 17865 8993 17877 8996
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 17954 8984 17960 9036
rect 18012 8984 18018 9036
rect 18230 8984 18236 9036
rect 18288 8984 18294 9036
rect 18414 8984 18420 9036
rect 18472 8984 18478 9036
rect 16114 8956 16120 8968
rect 15856 8928 16120 8956
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16666 8916 16672 8968
rect 16724 8916 16730 8968
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8925 17279 8959
rect 17221 8919 17279 8925
rect 9858 8888 9864 8900
rect 9508 8860 9864 8888
rect 9858 8848 9864 8860
rect 9916 8888 9922 8900
rect 12345 8891 12403 8897
rect 12345 8888 12357 8891
rect 9916 8860 12357 8888
rect 9916 8848 9922 8860
rect 12345 8857 12357 8860
rect 12391 8857 12403 8891
rect 12345 8851 12403 8857
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 13078 8888 13084 8900
rect 12492 8860 13084 8888
rect 12492 8848 12498 8860
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 14277 8891 14335 8897
rect 14277 8888 14289 8891
rect 13188 8860 14289 8888
rect 7926 8780 7932 8832
rect 7984 8780 7990 8832
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 13188 8820 13216 8860
rect 14277 8857 14289 8860
rect 14323 8857 14335 8891
rect 14277 8851 14335 8857
rect 16206 8848 16212 8900
rect 16264 8888 16270 8900
rect 17236 8888 17264 8919
rect 17954 8888 17960 8900
rect 16264 8860 17172 8888
rect 17236 8860 17960 8888
rect 16264 8848 16270 8860
rect 11848 8792 13216 8820
rect 11848 8780 11854 8792
rect 15286 8780 15292 8832
rect 15344 8820 15350 8832
rect 16022 8820 16028 8832
rect 15344 8792 16028 8820
rect 15344 8780 15350 8792
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16356 8792 17049 8820
rect 16356 8780 16362 8792
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 17144 8820 17172 8860
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 18233 8891 18291 8897
rect 18233 8888 18245 8891
rect 18012 8860 18245 8888
rect 18012 8848 18018 8860
rect 18233 8857 18245 8860
rect 18279 8857 18291 8891
rect 18233 8851 18291 8857
rect 18141 8823 18199 8829
rect 18141 8820 18153 8823
rect 17144 8792 18153 8820
rect 17037 8783 17095 8789
rect 18141 8789 18153 8792
rect 18187 8789 18199 8823
rect 18141 8783 18199 8789
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 11790 8576 11796 8628
rect 11848 8576 11854 8628
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 13170 8616 13176 8628
rect 12943 8588 13176 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 15381 8619 15439 8625
rect 15381 8616 15393 8619
rect 13872 8588 15393 8616
rect 13872 8576 13878 8588
rect 15381 8585 15393 8588
rect 15427 8585 15439 8619
rect 15381 8579 15439 8585
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16298 8616 16304 8628
rect 15988 8588 16304 8616
rect 15988 8576 15994 8588
rect 16298 8576 16304 8588
rect 16356 8576 16362 8628
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 16577 8619 16635 8625
rect 16577 8616 16589 8619
rect 16540 8588 16589 8616
rect 16540 8576 16546 8588
rect 16577 8585 16589 8588
rect 16623 8585 16635 8619
rect 16577 8579 16635 8585
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8548 8539 8551
rect 8570 8548 8576 8560
rect 8527 8520 8576 8548
rect 8527 8517 8539 8520
rect 8481 8511 8539 8517
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 12713 8551 12771 8557
rect 12713 8548 12725 8551
rect 11900 8520 12725 8548
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 11609 8483 11667 8489
rect 11609 8449 11621 8483
rect 11655 8480 11667 8483
rect 11698 8480 11704 8492
rect 11655 8452 11704 8480
rect 11655 8449 11667 8452
rect 11609 8443 11667 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 11900 8421 11928 8520
rect 12713 8517 12725 8520
rect 12759 8517 12771 8551
rect 12713 8511 12771 8517
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 14645 8551 14703 8557
rect 14645 8548 14657 8551
rect 14240 8520 14657 8548
rect 14240 8508 14246 8520
rect 14645 8517 14657 8520
rect 14691 8517 14703 8551
rect 16945 8551 17003 8557
rect 16945 8548 16957 8551
rect 14645 8511 14703 8517
rect 15028 8520 16957 8548
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 14734 8480 14740 8492
rect 14292 8452 14740 8480
rect 9594 8415 9652 8421
rect 9594 8412 9606 8415
rect 8904 8384 9606 8412
rect 8904 8372 8910 8384
rect 9594 8381 9606 8384
rect 9640 8381 9652 8415
rect 9594 8375 9652 8381
rect 11885 8415 11943 8421
rect 11885 8381 11897 8415
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 12158 8372 12164 8424
rect 12216 8372 12222 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12434 8412 12440 8424
rect 12299 8384 12440 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 10778 8304 10784 8356
rect 10836 8344 10842 8356
rect 11609 8347 11667 8353
rect 11609 8344 11621 8347
rect 10836 8316 11621 8344
rect 10836 8304 10842 8316
rect 11609 8313 11621 8316
rect 11655 8313 11667 8347
rect 12544 8344 12572 8440
rect 13541 8415 13599 8421
rect 13541 8412 13553 8415
rect 12912 8384 13553 8412
rect 12912 8353 12940 8384
rect 13541 8381 13553 8384
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13630 8372 13636 8424
rect 13688 8412 13694 8424
rect 14001 8415 14059 8421
rect 14001 8412 14013 8415
rect 13688 8384 14013 8412
rect 13688 8372 13694 8384
rect 14001 8381 14013 8384
rect 14047 8412 14059 8415
rect 14090 8412 14096 8424
rect 14047 8384 14096 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14292 8421 14320 8452
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 14277 8415 14335 8421
rect 14277 8381 14289 8415
rect 14323 8381 14335 8415
rect 14277 8375 14335 8381
rect 14369 8415 14427 8421
rect 14369 8381 14381 8415
rect 14415 8412 14427 8415
rect 14458 8412 14464 8424
rect 14415 8384 14464 8412
rect 14415 8381 14427 8384
rect 14369 8375 14427 8381
rect 12865 8347 12940 8353
rect 12865 8344 12877 8347
rect 12544 8316 12877 8344
rect 11609 8307 11667 8313
rect 12865 8313 12877 8316
rect 12911 8316 12940 8347
rect 12911 8313 12923 8316
rect 12865 8307 12923 8313
rect 13078 8304 13084 8356
rect 13136 8304 13142 8356
rect 13722 8304 13728 8356
rect 13780 8304 13786 8356
rect 13906 8304 13912 8356
rect 13964 8304 13970 8356
rect 14200 8344 14228 8375
rect 14458 8372 14464 8384
rect 14516 8412 14522 8424
rect 14516 8384 14872 8412
rect 14516 8372 14522 8384
rect 14737 8347 14795 8353
rect 14737 8344 14749 8347
rect 14200 8316 14749 8344
rect 14737 8313 14749 8316
rect 14783 8313 14795 8347
rect 14844 8344 14872 8384
rect 14918 8372 14924 8424
rect 14976 8372 14982 8424
rect 15028 8421 15056 8520
rect 16945 8517 16957 8520
rect 16991 8548 17003 8551
rect 17034 8548 17040 8560
rect 16991 8520 17040 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 17494 8508 17500 8560
rect 17552 8548 17558 8560
rect 17862 8548 17868 8560
rect 17552 8520 17868 8548
rect 17552 8508 17558 8520
rect 17862 8508 17868 8520
rect 17920 8548 17926 8560
rect 17920 8520 18184 8548
rect 17920 8508 17926 8520
rect 15838 8440 15844 8492
rect 15896 8480 15902 8492
rect 16669 8483 16727 8489
rect 15896 8452 16252 8480
rect 15896 8440 15902 8452
rect 15013 8415 15071 8421
rect 15013 8381 15025 8415
rect 15059 8381 15071 8415
rect 15013 8375 15071 8381
rect 15194 8372 15200 8424
rect 15252 8372 15258 8424
rect 15286 8372 15292 8424
rect 15344 8372 15350 8424
rect 15378 8372 15384 8424
rect 15436 8372 15442 8424
rect 15562 8372 15568 8424
rect 15620 8372 15626 8424
rect 15654 8372 15660 8424
rect 15712 8372 15718 8424
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8412 15991 8415
rect 16114 8412 16120 8424
rect 15979 8384 16120 8412
rect 15979 8381 15991 8384
rect 15933 8375 15991 8381
rect 15396 8344 15424 8372
rect 14844 8316 15424 8344
rect 14737 8307 14795 8313
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 15948 8344 15976 8375
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 15528 8316 15976 8344
rect 16224 8344 16252 8452
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 17770 8480 17776 8492
rect 16715 8452 17776 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 17770 8440 17776 8452
rect 17828 8480 17834 8492
rect 18156 8489 18184 8520
rect 18141 8483 18199 8489
rect 17828 8452 18000 8480
rect 17828 8440 17834 8452
rect 16574 8372 16580 8424
rect 16632 8372 16638 8424
rect 17221 8415 17279 8421
rect 17221 8381 17233 8415
rect 17267 8412 17279 8415
rect 17402 8412 17408 8424
rect 17267 8384 17408 8412
rect 17267 8381 17279 8384
rect 17221 8375 17279 8381
rect 17402 8372 17408 8384
rect 17460 8372 17466 8424
rect 17972 8421 18000 8452
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 17497 8415 17555 8421
rect 17497 8381 17509 8415
rect 17543 8381 17555 8415
rect 17497 8375 17555 8381
rect 17957 8415 18015 8421
rect 17957 8381 17969 8415
rect 18003 8412 18015 8415
rect 18414 8412 18420 8424
rect 18003 8384 18420 8412
rect 18003 8381 18015 8384
rect 17957 8375 18015 8381
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 16224 8316 17049 8344
rect 15528 8304 15534 8316
rect 17037 8313 17049 8316
rect 17083 8313 17095 8347
rect 17037 8307 17095 8313
rect 17310 8304 17316 8356
rect 17368 8344 17374 8356
rect 17512 8344 17540 8375
rect 18414 8372 18420 8384
rect 18472 8372 18478 8424
rect 17368 8316 18092 8344
rect 17368 8304 17374 8316
rect 11974 8236 11980 8288
rect 12032 8236 12038 8288
rect 12437 8279 12495 8285
rect 12437 8245 12449 8279
rect 12483 8276 12495 8279
rect 13262 8276 13268 8288
rect 12483 8248 13268 8276
rect 12483 8245 12495 8248
rect 12437 8239 12495 8245
rect 13262 8236 13268 8248
rect 13320 8236 13326 8288
rect 17405 8279 17463 8285
rect 17405 8245 17417 8279
rect 17451 8276 17463 8279
rect 17494 8276 17500 8288
rect 17451 8248 17500 8276
rect 17451 8245 17463 8248
rect 17405 8239 17463 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 17586 8236 17592 8288
rect 17644 8236 17650 8288
rect 18064 8285 18092 8316
rect 18049 8279 18107 8285
rect 18049 8245 18061 8279
rect 18095 8276 18107 8279
rect 18230 8276 18236 8288
rect 18095 8248 18236 8276
rect 18095 8245 18107 8248
rect 18049 8239 18107 8245
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 9953 8075 10011 8081
rect 9953 8041 9965 8075
rect 9999 8072 10011 8075
rect 10226 8072 10232 8084
rect 9999 8044 10232 8072
rect 9999 8041 10011 8044
rect 9953 8035 10011 8041
rect 10226 8032 10232 8044
rect 10284 8032 10290 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 11333 8075 11391 8081
rect 11333 8072 11345 8075
rect 10652 8044 11345 8072
rect 10652 8032 10658 8044
rect 11333 8041 11345 8044
rect 11379 8041 11391 8075
rect 11333 8035 11391 8041
rect 12158 8032 12164 8084
rect 12216 8032 12222 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13265 8075 13323 8081
rect 12492 8044 13124 8072
rect 12492 8032 12498 8044
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 9769 8007 9827 8013
rect 9769 8004 9781 8007
rect 9640 7976 9781 8004
rect 9640 7964 9646 7976
rect 9769 7973 9781 7976
rect 9815 7973 9827 8007
rect 9769 7967 9827 7973
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 10962 8004 10968 8016
rect 10376 7976 10968 8004
rect 10376 7964 10382 7976
rect 10962 7964 10968 7976
rect 11020 8004 11026 8016
rect 11425 8007 11483 8013
rect 11425 8004 11437 8007
rect 11020 7976 11437 8004
rect 11020 7964 11026 7976
rect 11425 7973 11437 7976
rect 11471 7973 11483 8007
rect 12897 8007 12955 8013
rect 12897 8004 12909 8007
rect 11425 7967 11483 7973
rect 12636 7976 12909 8004
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 12437 7939 12495 7945
rect 10091 7908 11008 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10980 7809 11008 7908
rect 12437 7905 12449 7939
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11974 7868 11980 7880
rect 11655 7840 11980 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 10965 7803 11023 7809
rect 10965 7769 10977 7803
rect 11011 7769 11023 7803
rect 12452 7800 12480 7899
rect 12526 7896 12532 7948
rect 12584 7896 12590 7948
rect 12636 7945 12664 7976
rect 12897 7973 12909 7976
rect 12943 7973 12955 8007
rect 12897 7967 12955 7973
rect 12621 7939 12679 7945
rect 12621 7905 12633 7939
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 12802 7896 12808 7948
rect 12860 7896 12866 7948
rect 13096 7945 13124 8044
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13354 8072 13360 8084
rect 13311 8044 13360 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13354 8032 13360 8044
rect 13412 8032 13418 8084
rect 14645 8075 14703 8081
rect 14645 8041 14657 8075
rect 14691 8072 14703 8075
rect 14918 8072 14924 8084
rect 14691 8044 14924 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 17865 8075 17923 8081
rect 17865 8072 17877 8075
rect 15712 8044 17877 8072
rect 15712 8032 15718 8044
rect 17865 8041 17877 8044
rect 17911 8041 17923 8075
rect 17865 8035 17923 8041
rect 13372 8004 13400 8032
rect 15194 8004 15200 8016
rect 13372 7976 15200 8004
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7936 13415 7939
rect 13446 7936 13452 7948
rect 13403 7908 13452 7936
rect 13403 7905 13415 7908
rect 13357 7899 13415 7905
rect 13096 7868 13124 7899
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13740 7945 13768 7976
rect 15194 7964 15200 7976
rect 15252 8004 15258 8016
rect 15289 8007 15347 8013
rect 15289 8004 15301 8007
rect 15252 7976 15301 8004
rect 15252 7964 15258 7976
rect 15289 7973 15301 7976
rect 15335 7973 15347 8007
rect 15289 7967 15347 7973
rect 15519 7973 15577 7979
rect 15519 7970 15531 7973
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7905 13783 7939
rect 13725 7899 13783 7905
rect 14458 7896 14464 7948
rect 14516 7896 14522 7948
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 13630 7868 13636 7880
rect 13096 7840 13636 7868
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 14660 7868 14688 7899
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15509 7939 15531 7970
rect 15565 7939 15577 7973
rect 17788 7976 18092 8004
rect 15509 7936 15577 7939
rect 14976 7933 15577 7936
rect 14976 7908 15537 7933
rect 14976 7896 14982 7908
rect 15304 7880 15332 7908
rect 17034 7896 17040 7948
rect 17092 7896 17098 7948
rect 17221 7939 17279 7945
rect 17221 7936 17233 7939
rect 17144 7908 17233 7936
rect 15010 7868 15016 7880
rect 14660 7840 15016 7868
rect 14660 7800 14688 7840
rect 15010 7828 15016 7840
rect 15068 7828 15074 7880
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 15930 7828 15936 7880
rect 15988 7868 15994 7880
rect 17144 7868 17172 7908
rect 17221 7905 17233 7908
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 17310 7896 17316 7948
rect 17368 7896 17374 7948
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7936 17463 7939
rect 17494 7936 17500 7948
rect 17451 7908 17500 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 17788 7945 17816 7976
rect 17773 7939 17831 7945
rect 17773 7936 17785 7939
rect 17644 7908 17785 7936
rect 17644 7896 17650 7908
rect 17773 7905 17785 7908
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 17954 7896 17960 7948
rect 18012 7896 18018 7948
rect 18064 7945 18092 7976
rect 18049 7939 18107 7945
rect 18049 7905 18061 7939
rect 18095 7905 18107 7939
rect 18049 7899 18107 7905
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7905 18291 7939
rect 18233 7899 18291 7905
rect 15988 7840 17172 7868
rect 15988 7828 15994 7840
rect 12452 7772 14688 7800
rect 17144 7800 17172 7840
rect 18248 7800 18276 7899
rect 17144 7772 18276 7800
rect 10965 7763 11023 7769
rect 9769 7735 9827 7741
rect 9769 7701 9781 7735
rect 9815 7732 9827 7735
rect 10226 7732 10232 7744
rect 9815 7704 10232 7732
rect 9815 7701 9827 7704
rect 9769 7695 9827 7701
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 13262 7692 13268 7744
rect 13320 7732 13326 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 13320 7704 13553 7732
rect 13320 7692 13326 7704
rect 13541 7701 13553 7704
rect 13587 7732 13599 7735
rect 13722 7732 13728 7744
rect 13587 7704 13728 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 15470 7692 15476 7744
rect 15528 7692 15534 7744
rect 15654 7692 15660 7744
rect 15712 7692 15718 7744
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 17681 7735 17739 7741
rect 17681 7732 17693 7735
rect 17552 7704 17693 7732
rect 17552 7692 17558 7704
rect 17681 7701 17693 7704
rect 17727 7701 17739 7735
rect 17681 7695 17739 7701
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 12802 7528 12808 7540
rect 12268 7500 12808 7528
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9732 7364 10057 7392
rect 9732 7352 9738 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 12268 7401 12296 7500
rect 12802 7488 12808 7500
rect 12860 7488 12866 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 17218 7528 17224 7540
rect 14332 7500 17224 7528
rect 14332 7488 14338 7500
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 18046 7528 18052 7540
rect 17451 7500 18052 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 15930 7460 15936 7472
rect 14292 7432 15936 7460
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 10652 7364 11069 7392
rect 10652 7352 10658 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 11287 7364 12265 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14292 7392 14320 7432
rect 15930 7420 15936 7432
rect 15988 7460 15994 7472
rect 15988 7432 16068 7460
rect 15988 7420 15994 7432
rect 15746 7392 15752 7404
rect 13872 7364 14320 7392
rect 13872 7352 13878 7364
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9088 7296 9781 7324
rect 9088 7284 9094 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 10962 7284 10968 7336
rect 11020 7284 11026 7336
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 11756 7296 12449 7324
rect 11756 7284 11762 7296
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 8386 7216 8392 7268
rect 8444 7216 8450 7268
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10560 7160 10609 7188
rect 10560 7148 10566 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 12452 7188 12480 7287
rect 12710 7284 12716 7336
rect 12768 7284 12774 7336
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7256 12679 7259
rect 13078 7256 13084 7268
rect 12667 7228 13084 7256
rect 12667 7225 12679 7228
rect 12621 7219 12679 7225
rect 13078 7216 13084 7228
rect 13136 7256 13142 7268
rect 13924 7256 13952 7287
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14292 7333 14320 7364
rect 14936 7364 15752 7392
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 14056 7296 14105 7324
rect 14056 7284 14062 7296
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14200 7256 14228 7287
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 14936 7324 14964 7364
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 14516 7296 14964 7324
rect 14516 7284 14522 7296
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15838 7324 15844 7336
rect 15068 7296 15844 7324
rect 15068 7284 15074 7296
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16040 7333 16068 7432
rect 17494 7352 17500 7404
rect 17552 7352 17558 7404
rect 16025 7327 16083 7333
rect 16025 7293 16037 7327
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16574 7324 16580 7336
rect 16347 7296 16580 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 14369 7259 14427 7265
rect 14369 7256 14381 7259
rect 13136 7228 14136 7256
rect 14200 7228 14381 7256
rect 13136 7216 13142 7228
rect 13170 7188 13176 7200
rect 12452 7160 13176 7188
rect 10597 7151 10655 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13725 7191 13783 7197
rect 13725 7157 13737 7191
rect 13771 7188 13783 7191
rect 13998 7188 14004 7200
rect 13771 7160 14004 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 13998 7148 14004 7160
rect 14056 7148 14062 7200
rect 14108 7188 14136 7228
rect 14369 7225 14381 7228
rect 14415 7225 14427 7259
rect 14369 7219 14427 7225
rect 15102 7216 15108 7268
rect 15160 7256 15166 7268
rect 15197 7259 15255 7265
rect 15197 7256 15209 7259
rect 15160 7228 15209 7256
rect 15160 7216 15166 7228
rect 15197 7225 15209 7228
rect 15243 7225 15255 7259
rect 15197 7219 15255 7225
rect 15286 7216 15292 7268
rect 15344 7256 15350 7268
rect 17037 7259 17095 7265
rect 17037 7256 17049 7259
rect 15344 7228 17049 7256
rect 15344 7216 15350 7228
rect 17037 7225 17049 7228
rect 17083 7225 17095 7259
rect 17037 7219 17095 7225
rect 14274 7188 14280 7200
rect 14108 7160 14280 7188
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 15381 7191 15439 7197
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15470 7188 15476 7200
rect 15427 7160 15476 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 15838 7188 15844 7200
rect 15620 7160 15844 7188
rect 15620 7148 15626 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16209 7191 16267 7197
rect 16209 7157 16221 7191
rect 16255 7188 16267 7191
rect 16850 7188 16856 7200
rect 16255 7160 16856 7188
rect 16255 7157 16267 7160
rect 16209 7151 16267 7157
rect 16850 7148 16856 7160
rect 16908 7188 16914 7200
rect 17402 7188 17408 7200
rect 16908 7160 17408 7188
rect 16908 7148 16914 7160
rect 17402 7148 17408 7160
rect 17460 7148 17466 7200
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 10045 6987 10103 6993
rect 10045 6953 10057 6987
rect 10091 6984 10103 6987
rect 10134 6984 10140 6996
rect 10091 6956 10140 6984
rect 10091 6953 10103 6956
rect 10045 6947 10103 6953
rect 10134 6944 10140 6956
rect 10192 6984 10198 6996
rect 10594 6984 10600 6996
rect 10192 6956 10600 6984
rect 10192 6944 10198 6956
rect 10594 6944 10600 6956
rect 10652 6984 10658 6996
rect 11425 6987 11483 6993
rect 11425 6984 11437 6987
rect 10652 6956 11437 6984
rect 10652 6944 10658 6956
rect 11425 6953 11437 6956
rect 11471 6953 11483 6987
rect 11425 6947 11483 6953
rect 13170 6944 13176 6996
rect 13228 6984 13234 6996
rect 13538 6984 13544 6996
rect 13228 6956 13544 6984
rect 13228 6944 13234 6956
rect 13538 6944 13544 6956
rect 13596 6984 13602 6996
rect 13596 6956 13952 6984
rect 13596 6944 13602 6956
rect 8864 6888 9536 6916
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8864 6848 8892 6888
rect 8803 6820 8892 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 9232 6848 9260 6888
rect 9171 6820 9260 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 9048 6780 9076 6811
rect 9306 6808 9312 6860
rect 9364 6808 9370 6860
rect 9398 6808 9404 6860
rect 9456 6808 9462 6860
rect 9508 6848 9536 6888
rect 9950 6876 9956 6928
rect 10008 6916 10014 6928
rect 10962 6916 10968 6928
rect 10008 6888 10968 6916
rect 10008 6876 10014 6888
rect 10962 6876 10968 6888
rect 11020 6916 11026 6928
rect 11333 6919 11391 6925
rect 11333 6916 11345 6919
rect 11020 6888 11345 6916
rect 11020 6876 11026 6888
rect 11333 6885 11345 6888
rect 11379 6885 11391 6919
rect 11333 6879 11391 6885
rect 13265 6919 13323 6925
rect 13265 6885 13277 6919
rect 13311 6916 13323 6919
rect 13446 6916 13452 6928
rect 13311 6888 13452 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 13924 6916 13952 6956
rect 14642 6944 14648 6996
rect 14700 6944 14706 6996
rect 14752 6956 15700 6984
rect 14752 6916 14780 6956
rect 13924 6888 14780 6916
rect 9582 6848 9588 6860
rect 9508 6820 9588 6848
rect 9582 6808 9588 6820
rect 9640 6848 9646 6860
rect 9640 6820 10180 6848
rect 9640 6808 9646 6820
rect 9048 6752 9628 6780
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9030 6712 9036 6724
rect 8803 6684 9036 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9030 6672 9036 6684
rect 9088 6672 9094 6724
rect 9600 6721 9628 6752
rect 9585 6715 9643 6721
rect 9585 6681 9597 6715
rect 9631 6681 9643 6715
rect 10152 6712 10180 6820
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10686 6848 10692 6860
rect 10643 6820 10692 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 10778 6808 10784 6860
rect 10836 6808 10842 6860
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 12345 6851 12403 6857
rect 12345 6817 12357 6851
rect 12391 6848 12403 6851
rect 12618 6848 12624 6860
rect 12391 6820 12624 6848
rect 12391 6817 12403 6820
rect 12345 6811 12403 6817
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12768 6820 12909 6848
rect 12768 6808 12774 6820
rect 12897 6817 12909 6820
rect 12943 6848 12955 6851
rect 12943 6820 13676 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6780 10287 6783
rect 11146 6780 11152 6792
rect 10275 6752 11152 6780
rect 10275 6749 10287 6752
rect 10229 6743 10287 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 11609 6783 11667 6789
rect 11609 6749 11621 6783
rect 11655 6780 11667 6783
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11655 6752 11989 6780
rect 11655 6749 11667 6752
rect 11609 6743 11667 6749
rect 11977 6749 11989 6752
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12253 6783 12311 6789
rect 12253 6749 12265 6783
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12805 6783 12863 6789
rect 12483 6752 12664 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 10686 6712 10692 6724
rect 10152 6684 10692 6712
rect 9585 6675 9643 6681
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 11238 6712 11244 6724
rect 10827 6684 11244 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 12268 6712 12296 6743
rect 12526 6712 12532 6724
rect 12268 6684 12532 6712
rect 12526 6672 12532 6684
rect 12584 6672 12590 6724
rect 12636 6721 12664 6752
rect 12805 6749 12817 6783
rect 12851 6749 12863 6783
rect 12805 6743 12863 6749
rect 12621 6715 12679 6721
rect 12621 6681 12633 6715
rect 12667 6681 12679 6715
rect 12621 6675 12679 6681
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 12820 6712 12848 6743
rect 13170 6740 13176 6792
rect 13228 6740 13234 6792
rect 13648 6780 13676 6820
rect 13722 6808 13728 6860
rect 13780 6808 13786 6860
rect 14016 6857 14044 6888
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6817 14059 6851
rect 14001 6811 14059 6817
rect 14366 6808 14372 6860
rect 14424 6808 14430 6860
rect 14642 6851 14700 6857
rect 14642 6817 14654 6851
rect 14688 6848 14700 6851
rect 14752 6848 14780 6888
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15436 6888 15608 6916
rect 15436 6876 15442 6888
rect 14688 6820 14780 6848
rect 15105 6851 15163 6857
rect 14688 6817 14700 6820
rect 14642 6811 14700 6817
rect 15105 6817 15117 6851
rect 15151 6848 15163 6851
rect 15286 6848 15292 6860
rect 15151 6820 15292 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 15286 6808 15292 6820
rect 15344 6808 15350 6860
rect 15470 6808 15476 6860
rect 15528 6808 15534 6860
rect 15580 6857 15608 6888
rect 15672 6857 15700 6956
rect 16022 6944 16028 6996
rect 16080 6984 16086 6996
rect 16869 6987 16927 6993
rect 16869 6984 16881 6987
rect 16080 6956 16881 6984
rect 16080 6944 16086 6956
rect 16869 6953 16881 6956
rect 16915 6953 16927 6987
rect 16869 6947 16927 6953
rect 16666 6876 16672 6928
rect 16724 6876 16730 6928
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 13817 6783 13875 6789
rect 13817 6780 13829 6783
rect 13648 6752 13829 6780
rect 13817 6749 13829 6752
rect 13863 6780 13875 6783
rect 15010 6780 15016 6792
rect 13863 6752 15016 6780
rect 13863 6749 13875 6752
rect 13817 6743 13875 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 15252 6752 15393 6780
rect 15252 6740 15258 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 13909 6715 13967 6721
rect 12768 6684 13768 6712
rect 12768 6672 12774 6684
rect 13740 6656 13768 6684
rect 13909 6681 13921 6715
rect 13955 6712 13967 6715
rect 14277 6715 14335 6721
rect 14277 6712 14289 6715
rect 13955 6684 14289 6712
rect 13955 6681 13967 6684
rect 13909 6675 13967 6681
rect 14277 6681 14289 6684
rect 14323 6681 14335 6715
rect 15580 6712 15608 6811
rect 14277 6675 14335 6681
rect 14384 6684 15608 6712
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9490 6644 9496 6656
rect 9171 6616 9496 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 10962 6604 10968 6656
rect 11020 6604 11026 6656
rect 13538 6604 13544 6656
rect 13596 6604 13602 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 14384 6644 14412 6684
rect 13780 6616 14412 6644
rect 13780 6604 13786 6616
rect 14458 6604 14464 6656
rect 14516 6604 14522 6656
rect 15013 6647 15071 6653
rect 15013 6613 15025 6647
rect 15059 6644 15071 6647
rect 15197 6647 15255 6653
rect 15197 6644 15209 6647
rect 15059 6616 15209 6644
rect 15059 6613 15071 6616
rect 15013 6607 15071 6613
rect 15197 6613 15209 6616
rect 15243 6613 15255 6647
rect 15197 6607 15255 6613
rect 16850 6604 16856 6656
rect 16908 6604 16914 6656
rect 17037 6647 17095 6653
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17310 6644 17316 6656
rect 17083 6616 17316 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9456 6412 9689 6440
rect 9456 6400 9462 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 9677 6403 9735 6409
rect 10336 6412 14381 6440
rect 10134 6264 10140 6316
rect 10192 6264 10198 6316
rect 10336 6313 10364 6412
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14700 6412 15117 6440
rect 14700 6400 14706 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15838 6440 15844 6452
rect 15105 6403 15163 6409
rect 15304 6412 15844 6440
rect 11054 6332 11060 6384
rect 11112 6332 11118 6384
rect 11146 6332 11152 6384
rect 11204 6372 11210 6384
rect 14458 6372 14464 6384
rect 11204 6344 14464 6372
rect 11204 6332 11210 6344
rect 14458 6332 14464 6344
rect 14516 6332 14522 6384
rect 14921 6375 14979 6381
rect 14921 6341 14933 6375
rect 14967 6372 14979 6375
rect 15194 6372 15200 6384
rect 14967 6344 15200 6372
rect 14967 6341 14979 6344
rect 14921 6335 14979 6341
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 10321 6307 10379 6313
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10744 6276 11100 6304
rect 10744 6264 10750 6276
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10045 6239 10103 6245
rect 10045 6236 10057 6239
rect 10008 6208 10057 6236
rect 10008 6196 10014 6208
rect 10045 6205 10057 6208
rect 10091 6205 10103 6239
rect 10045 6199 10103 6205
rect 10781 6239 10839 6245
rect 10781 6205 10793 6239
rect 10827 6236 10839 6239
rect 10962 6236 10968 6248
rect 10827 6208 10968 6236
rect 10827 6205 10839 6208
rect 10781 6199 10839 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11072 6245 11100 6276
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 15304 6313 15332 6412
rect 15838 6400 15844 6412
rect 15896 6400 15902 6452
rect 16945 6443 17003 6449
rect 16945 6409 16957 6443
rect 16991 6440 17003 6443
rect 17310 6440 17316 6452
rect 16991 6412 17316 6440
rect 16991 6409 17003 6412
rect 16945 6403 17003 6409
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 15470 6372 15476 6384
rect 15396 6344 15476 6372
rect 15396 6313 15424 6344
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 16761 6375 16819 6381
rect 16761 6341 16773 6375
rect 16807 6341 16819 6375
rect 17221 6375 17279 6381
rect 17221 6372 17233 6375
rect 16761 6335 16819 6341
rect 17144 6344 17233 6372
rect 15289 6307 15347 6313
rect 12584 6276 14872 6304
rect 12584 6264 12590 6276
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 13538 6196 13544 6248
rect 13596 6236 13602 6248
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13596 6208 13829 6236
rect 13596 6196 13602 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13998 6196 14004 6248
rect 14056 6196 14062 6248
rect 14182 6196 14188 6248
rect 14240 6196 14246 6248
rect 14844 6245 14872 6276
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 15654 6304 15660 6316
rect 15611 6276 15660 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 15804 6276 16313 6304
rect 15804 6264 15810 6276
rect 16301 6273 16313 6276
rect 16347 6273 16359 6307
rect 16301 6267 16359 6273
rect 14829 6239 14887 6245
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 14918 6236 14924 6248
rect 14875 6208 14924 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6236 15071 6239
rect 15102 6236 15108 6248
rect 15059 6208 15108 6236
rect 15059 6205 15071 6208
rect 15013 6199 15071 6205
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6236 15531 6239
rect 16393 6239 16451 6245
rect 15519 6208 15700 6236
rect 15519 6205 15531 6208
rect 15473 6199 15531 6205
rect 10870 6128 10876 6180
rect 10928 6128 10934 6180
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6168 14151 6171
rect 15672 6168 15700 6208
rect 16393 6205 16405 6239
rect 16439 6236 16451 6239
rect 16574 6236 16580 6248
rect 16439 6208 16580 6236
rect 16439 6205 16451 6208
rect 16393 6199 16451 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16776 6236 16804 6335
rect 17144 6313 17172 6344
rect 17221 6341 17233 6344
rect 17267 6341 17279 6375
rect 17221 6335 17279 6341
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 16853 6239 16911 6245
rect 16853 6236 16865 6239
rect 16776 6208 16865 6236
rect 16853 6205 16865 6208
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 16758 6168 16764 6180
rect 14139 6140 15608 6168
rect 15672 6140 16764 6168
rect 14139 6137 14151 6140
rect 14093 6131 14151 6137
rect 15580 6100 15608 6140
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 16868 6168 16896 6199
rect 16942 6196 16948 6248
rect 17000 6236 17006 6248
rect 17218 6236 17224 6248
rect 17000 6208 17224 6236
rect 17000 6196 17006 6208
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 17310 6196 17316 6248
rect 17368 6236 17374 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 17368 6208 17509 6236
rect 17368 6196 17374 6208
rect 17497 6205 17509 6208
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 16868 6140 17448 6168
rect 17420 6109 17448 6140
rect 17129 6103 17187 6109
rect 17129 6100 17141 6103
rect 15580 6072 17141 6100
rect 17129 6069 17141 6072
rect 17175 6069 17187 6103
rect 17129 6063 17187 6069
rect 17405 6103 17463 6109
rect 17405 6069 17417 6103
rect 17451 6069 17463 6103
rect 17405 6063 17463 6069
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9732 5800 10088 5828
rect 9732 5788 9738 5800
rect 9490 5720 9496 5772
rect 9548 5760 9554 5772
rect 10060 5769 10088 5800
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11578 5831 11636 5837
rect 11578 5828 11590 5831
rect 11112 5800 11590 5828
rect 11112 5788 11118 5800
rect 11578 5797 11590 5800
rect 11624 5797 11636 5831
rect 11578 5791 11636 5797
rect 9778 5763 9836 5769
rect 9778 5760 9790 5763
rect 9548 5732 9790 5760
rect 9548 5720 9554 5732
rect 9778 5729 9790 5732
rect 9824 5729 9836 5763
rect 9778 5723 9836 5729
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10962 5760 10968 5772
rect 10091 5732 10968 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 10962 5720 10968 5732
rect 11020 5760 11026 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11020 5732 11345 5760
rect 11020 5720 11026 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 13630 5556 13636 5568
rect 12759 5528 13636 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 9674 5352 9680 5364
rect 9416 5324 9680 5352
rect 9416 5225 9444 5324
rect 9674 5312 9680 5324
rect 9732 5312 9738 5364
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5185 9459 5219
rect 9401 5179 9459 5185
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 9668 5151 9726 5157
rect 9668 5117 9680 5151
rect 9714 5148 9726 5151
rect 10226 5148 10232 5160
rect 9714 5120 10232 5148
rect 9714 5117 9726 5120
rect 9668 5111 9726 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10980 5148 11008 5176
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 10980 5120 16681 5148
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 16669 5111 16727 5117
rect 11238 5089 11244 5092
rect 11232 5080 11244 5089
rect 11199 5052 11244 5080
rect 11232 5043 11244 5052
rect 11238 5040 11244 5043
rect 11296 5040 11302 5092
rect 11606 5040 11612 5092
rect 11664 5080 11670 5092
rect 16914 5083 16972 5089
rect 16914 5080 16926 5083
rect 11664 5052 16926 5080
rect 11664 5040 11670 5052
rect 16914 5049 16926 5052
rect 16960 5049 16972 5083
rect 16914 5043 16972 5049
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 11054 5012 11060 5024
rect 10827 4984 11060 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 12345 5015 12403 5021
rect 12345 4981 12357 5015
rect 12391 5012 12403 5015
rect 16114 5012 16120 5024
rect 12391 4984 16120 5012
rect 12391 4981 12403 4984
rect 12345 4975 12403 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 18049 5015 18107 5021
rect 18049 4981 18061 5015
rect 18095 5012 18107 5015
rect 18598 5012 18604 5024
rect 18095 4984 18604 5012
rect 18095 4981 18107 4984
rect 18049 4975 18107 4981
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 7926 4128 7932 4140
rect 3752 4100 7932 4128
rect 3752 4088 3758 4100
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 8662 3720 8668 3732
rect 6236 3692 8668 3720
rect 6236 3680 6242 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 1210 3612 1216 3664
rect 1268 3652 1274 3664
rect 8386 3652 8392 3664
rect 1268 3624 8392 3652
rect 1268 3612 1274 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 10508 18912 10560 18964
rect 848 18776 900 18828
rect 2504 18776 2556 18828
rect 4160 18776 4212 18828
rect 5816 18776 5868 18828
rect 7472 18776 7524 18828
rect 9128 18776 9180 18828
rect 11060 18776 11112 18828
rect 12440 18776 12492 18828
rect 14096 18776 14148 18828
rect 15752 18776 15804 18828
rect 17408 18776 17460 18828
rect 7196 18708 7248 18760
rect 8024 18640 8076 18692
rect 6920 18572 6972 18624
rect 8668 18572 8720 18624
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 10232 18572 10284 18624
rect 12624 18572 12676 18624
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 15200 18572 15252 18624
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 7012 18368 7064 18420
rect 10416 18300 10468 18352
rect 4160 18164 4212 18216
rect 7288 18164 7340 18216
rect 7564 18207 7616 18216
rect 7564 18173 7573 18207
rect 7573 18173 7607 18207
rect 7607 18173 7616 18207
rect 7564 18164 7616 18173
rect 5724 18071 5776 18080
rect 5724 18037 5733 18071
rect 5733 18037 5767 18071
rect 5767 18037 5776 18071
rect 5724 18028 5776 18037
rect 6276 18028 6328 18080
rect 7472 18096 7524 18148
rect 7104 18028 7156 18080
rect 7288 18071 7340 18080
rect 7288 18037 7297 18071
rect 7297 18037 7331 18071
rect 7331 18037 7340 18071
rect 7288 18028 7340 18037
rect 7380 18028 7432 18080
rect 9128 18164 9180 18216
rect 9680 18164 9732 18216
rect 10232 18207 10284 18216
rect 10232 18173 10241 18207
rect 10241 18173 10275 18207
rect 10275 18173 10284 18207
rect 10232 18164 10284 18173
rect 10508 18164 10560 18216
rect 17500 18164 17552 18216
rect 8852 18096 8904 18148
rect 7748 18028 7800 18080
rect 9680 18028 9732 18080
rect 10232 18071 10284 18080
rect 10232 18037 10241 18071
rect 10241 18037 10275 18071
rect 10275 18037 10284 18071
rect 10232 18028 10284 18037
rect 15844 18071 15896 18080
rect 15844 18037 15853 18071
rect 15853 18037 15887 18071
rect 15887 18037 15896 18071
rect 15844 18028 15896 18037
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 7380 17824 7432 17876
rect 7472 17824 7524 17876
rect 8852 17867 8904 17876
rect 8852 17833 8861 17867
rect 8861 17833 8895 17867
rect 8895 17833 8904 17867
rect 8852 17824 8904 17833
rect 4160 17688 4212 17740
rect 4344 17731 4396 17740
rect 4344 17697 4378 17731
rect 4378 17697 4396 17731
rect 4344 17688 4396 17697
rect 7196 17688 7248 17740
rect 10416 17756 10468 17808
rect 15844 17756 15896 17808
rect 16948 17756 17000 17808
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 8576 17731 8628 17740
rect 8576 17697 8585 17731
rect 8585 17697 8619 17731
rect 8619 17697 8628 17731
rect 8576 17688 8628 17697
rect 8668 17731 8720 17740
rect 8668 17697 8677 17731
rect 8677 17697 8711 17731
rect 8711 17697 8720 17731
rect 8668 17688 8720 17697
rect 8944 17731 8996 17740
rect 8944 17697 8953 17731
rect 8953 17697 8987 17731
rect 8987 17697 8996 17731
rect 8944 17688 8996 17697
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 7472 17663 7524 17672
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 7564 17620 7616 17672
rect 9496 17688 9548 17740
rect 10140 17688 10192 17740
rect 9128 17620 9180 17672
rect 5448 17595 5500 17604
rect 5448 17561 5457 17595
rect 5457 17561 5491 17595
rect 5491 17561 5500 17595
rect 5448 17552 5500 17561
rect 6920 17552 6972 17604
rect 7748 17552 7800 17604
rect 8944 17552 8996 17604
rect 15292 17620 15344 17672
rect 5816 17527 5868 17536
rect 5816 17493 5825 17527
rect 5825 17493 5859 17527
rect 5859 17493 5868 17527
rect 5816 17484 5868 17493
rect 7196 17484 7248 17536
rect 7472 17484 7524 17536
rect 7840 17484 7892 17536
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 8392 17484 8444 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 4344 17280 4396 17332
rect 7104 17280 7156 17332
rect 7932 17280 7984 17332
rect 8944 17280 8996 17332
rect 11336 17323 11388 17332
rect 11336 17289 11345 17323
rect 11345 17289 11379 17323
rect 11379 17289 11388 17323
rect 11336 17280 11388 17289
rect 7012 17212 7064 17264
rect 4252 17144 4304 17196
rect 5724 17144 5776 17196
rect 8576 17212 8628 17264
rect 1860 17076 1912 17128
rect 3700 17076 3752 17128
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 5816 17076 5868 17128
rect 7288 17144 7340 17196
rect 9312 17144 9364 17196
rect 9588 17144 9640 17196
rect 10416 17212 10468 17264
rect 10324 17144 10376 17196
rect 6276 17119 6328 17128
rect 6276 17085 6285 17119
rect 6285 17085 6319 17119
rect 6319 17085 6328 17119
rect 6276 17076 6328 17085
rect 7380 17076 7432 17128
rect 9680 17076 9732 17128
rect 10140 17119 10192 17128
rect 10140 17085 10149 17119
rect 10149 17085 10183 17119
rect 10183 17085 10192 17119
rect 10140 17076 10192 17085
rect 8668 17008 8720 17060
rect 10416 17119 10468 17128
rect 10416 17085 10425 17119
rect 10425 17085 10459 17119
rect 10459 17085 10468 17119
rect 10416 17076 10468 17085
rect 10692 17008 10744 17060
rect 16764 17008 16816 17060
rect 17868 17008 17920 17060
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 7196 16940 7248 16992
rect 10324 16983 10376 16992
rect 10324 16949 10333 16983
rect 10333 16949 10367 16983
rect 10367 16949 10376 16983
rect 10324 16940 10376 16949
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 4160 16736 4212 16788
rect 9680 16736 9732 16788
rect 2412 16668 2464 16720
rect 3700 16711 3752 16720
rect 3700 16677 3709 16711
rect 3709 16677 3743 16711
rect 3743 16677 3752 16711
rect 3700 16668 3752 16677
rect 7380 16668 7432 16720
rect 8024 16668 8076 16720
rect 11244 16668 11296 16720
rect 3976 16643 4028 16652
rect 3976 16609 3985 16643
rect 3985 16609 4019 16643
rect 4019 16609 4028 16643
rect 3976 16600 4028 16609
rect 4160 16643 4212 16652
rect 4160 16609 4169 16643
rect 4169 16609 4203 16643
rect 4203 16609 4212 16643
rect 4160 16600 4212 16609
rect 4436 16643 4488 16652
rect 4436 16609 4470 16643
rect 4470 16609 4488 16643
rect 4436 16600 4488 16609
rect 9496 16600 9548 16652
rect 10048 16643 10100 16652
rect 10048 16609 10057 16643
rect 10057 16609 10091 16643
rect 10091 16609 10100 16643
rect 10048 16600 10100 16609
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 3608 16464 3660 16516
rect 4160 16464 4212 16516
rect 5724 16532 5776 16584
rect 3516 16396 3568 16448
rect 3884 16439 3936 16448
rect 3884 16405 3893 16439
rect 3893 16405 3927 16439
rect 3927 16405 3936 16439
rect 3884 16396 3936 16405
rect 5816 16439 5868 16448
rect 5816 16405 5825 16439
rect 5825 16405 5859 16439
rect 5859 16405 5868 16439
rect 5816 16396 5868 16405
rect 7012 16396 7064 16448
rect 8208 16396 8260 16448
rect 10692 16396 10744 16448
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 3976 16192 4028 16244
rect 5448 16192 5500 16244
rect 3516 16124 3568 16176
rect 4620 16124 4672 16176
rect 2872 16056 2924 16108
rect 1860 16031 1912 16040
rect 1860 15997 1869 16031
rect 1869 15997 1903 16031
rect 1903 15997 1912 16031
rect 1860 15988 1912 15997
rect 2780 15988 2832 16040
rect 3516 15988 3568 16040
rect 3608 16031 3660 16040
rect 3608 15997 3617 16031
rect 3617 15997 3651 16031
rect 3651 15997 3660 16031
rect 5448 16056 5500 16108
rect 10048 16192 10100 16244
rect 11336 16192 11388 16244
rect 12532 16192 12584 16244
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 7932 16124 7984 16176
rect 12440 16124 12492 16176
rect 7012 16056 7064 16108
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 3608 15988 3660 15997
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2320 15852 2372 15904
rect 2596 15895 2648 15904
rect 2596 15861 2605 15895
rect 2605 15861 2639 15895
rect 2639 15861 2648 15895
rect 2596 15852 2648 15861
rect 2964 15920 3016 15972
rect 3332 15852 3384 15904
rect 5724 16031 5776 16040
rect 5724 15997 5733 16031
rect 5733 15997 5767 16031
rect 5767 15997 5776 16031
rect 5724 15988 5776 15997
rect 6460 15988 6512 16040
rect 6644 15920 6696 15972
rect 7380 16031 7432 16040
rect 7380 15997 7389 16031
rect 7389 15997 7423 16031
rect 7423 15997 7432 16031
rect 7380 15988 7432 15997
rect 13084 16056 13136 16108
rect 8116 15988 8168 16040
rect 9128 16031 9180 16040
rect 9128 15997 9137 16031
rect 9137 15997 9171 16031
rect 9171 15997 9180 16031
rect 9128 15988 9180 15997
rect 11060 16031 11112 16040
rect 11060 15997 11069 16031
rect 11069 15997 11103 16031
rect 11103 15997 11112 16031
rect 11060 15988 11112 15997
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 13268 15988 13320 16040
rect 14372 16031 14424 16040
rect 14372 15997 14381 16031
rect 14381 15997 14415 16031
rect 14415 15997 14424 16031
rect 14372 15988 14424 15997
rect 14924 15988 14976 16040
rect 8392 15920 8444 15972
rect 9220 15920 9272 15972
rect 12900 15920 12952 15972
rect 13452 15920 13504 15972
rect 7196 15852 7248 15904
rect 11980 15852 12032 15904
rect 12348 15852 12400 15904
rect 12808 15852 12860 15904
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 13544 15852 13596 15904
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 4436 15648 4488 15700
rect 6920 15648 6972 15700
rect 7380 15648 7432 15700
rect 7472 15648 7524 15700
rect 9220 15691 9272 15700
rect 9220 15657 9229 15691
rect 9229 15657 9263 15691
rect 9263 15657 9272 15691
rect 9220 15648 9272 15657
rect 9680 15648 9732 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 12808 15691 12860 15700
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 13636 15648 13688 15700
rect 15292 15648 15344 15700
rect 1676 15580 1728 15632
rect 2136 15512 2188 15564
rect 2596 15512 2648 15564
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 2780 15487 2832 15496
rect 2780 15453 2789 15487
rect 2789 15453 2823 15487
rect 2823 15453 2832 15487
rect 2780 15444 2832 15453
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 2872 15444 2924 15453
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3148 15444 3200 15496
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 4620 15512 4672 15564
rect 6736 15512 6788 15564
rect 7288 15580 7340 15632
rect 11704 15580 11756 15632
rect 5816 15444 5868 15496
rect 7104 15512 7156 15564
rect 8208 15555 8260 15564
rect 8208 15521 8217 15555
rect 8217 15521 8251 15555
rect 8251 15521 8260 15555
rect 8208 15512 8260 15521
rect 8300 15555 8352 15564
rect 8300 15521 8309 15555
rect 8309 15521 8343 15555
rect 8343 15521 8352 15555
rect 8300 15512 8352 15521
rect 8392 15555 8444 15564
rect 8392 15521 8401 15555
rect 8401 15521 8435 15555
rect 8435 15521 8444 15555
rect 8392 15512 8444 15521
rect 8944 15512 8996 15564
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 9588 15512 9640 15564
rect 3240 15376 3292 15428
rect 7840 15444 7892 15496
rect 2412 15308 2464 15360
rect 5448 15308 5500 15360
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 9496 15376 9548 15428
rect 8024 15308 8076 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 12440 15555 12492 15564
rect 12440 15521 12449 15555
rect 12449 15521 12483 15555
rect 12483 15521 12492 15555
rect 12440 15512 12492 15521
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 13360 15580 13412 15632
rect 11704 15376 11756 15428
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 13084 15308 13136 15360
rect 13268 15487 13320 15496
rect 13268 15453 13277 15487
rect 13277 15453 13311 15487
rect 13311 15453 13320 15487
rect 13268 15444 13320 15453
rect 13636 15555 13688 15564
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 13912 15555 13964 15564
rect 13912 15521 13946 15555
rect 13946 15521 13964 15555
rect 13912 15512 13964 15521
rect 13452 15444 13504 15496
rect 13452 15308 13504 15360
rect 13636 15308 13688 15360
rect 15108 15308 15160 15360
rect 15384 15351 15436 15360
rect 15384 15317 15393 15351
rect 15393 15317 15427 15351
rect 15427 15317 15436 15351
rect 15384 15308 15436 15317
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 2320 15104 2372 15156
rect 3148 15104 3200 15156
rect 3516 15104 3568 15156
rect 6184 15104 6236 15156
rect 1676 15036 1728 15088
rect 2320 14968 2372 15020
rect 4160 14968 4212 15020
rect 6368 14900 6420 14952
rect 9128 14900 9180 14952
rect 10692 14943 10744 14952
rect 10692 14909 10701 14943
rect 10701 14909 10735 14943
rect 10735 14909 10744 14943
rect 10692 14900 10744 14909
rect 11796 15104 11848 15156
rect 13176 15104 13228 15156
rect 11980 14968 12032 15020
rect 13084 15011 13136 15020
rect 13084 14977 13093 15011
rect 13093 14977 13127 15011
rect 13127 14977 13136 15011
rect 13084 14968 13136 14977
rect 14924 15104 14976 15156
rect 15108 15104 15160 15156
rect 16856 15147 16908 15156
rect 16856 15113 16865 15147
rect 16865 15113 16899 15147
rect 16899 15113 16908 15147
rect 16856 15104 16908 15113
rect 13452 15036 13504 15088
rect 14464 15036 14516 15088
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 12992 14943 13044 14952
rect 11704 14900 11756 14909
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 2412 14875 2464 14884
rect 2412 14841 2421 14875
rect 2421 14841 2455 14875
rect 2455 14841 2464 14875
rect 2412 14832 2464 14841
rect 3240 14832 3292 14884
rect 6184 14832 6236 14884
rect 7104 14832 7156 14884
rect 9496 14832 9548 14884
rect 11520 14832 11572 14884
rect 12900 14832 12952 14884
rect 13636 14900 13688 14952
rect 15292 14968 15344 15020
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 14096 14900 14148 14952
rect 16764 14900 16816 14952
rect 16948 14943 17000 14952
rect 16948 14909 16957 14943
rect 16957 14909 16991 14943
rect 16991 14909 17000 14943
rect 16948 14900 17000 14909
rect 14372 14832 14424 14884
rect 2136 14764 2188 14816
rect 3332 14764 3384 14816
rect 8116 14764 8168 14816
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 14924 14764 14976 14816
rect 17408 14832 17460 14884
rect 17132 14764 17184 14816
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 2044 14424 2096 14476
rect 2228 14467 2280 14476
rect 2228 14433 2262 14467
rect 2262 14433 2280 14467
rect 2228 14424 2280 14433
rect 4068 14424 4120 14476
rect 6184 14535 6236 14544
rect 6184 14501 6193 14535
rect 6193 14501 6227 14535
rect 6227 14501 6236 14535
rect 6184 14492 6236 14501
rect 4436 14467 4488 14476
rect 4436 14433 4445 14467
rect 4445 14433 4479 14467
rect 4479 14433 4488 14467
rect 4436 14424 4488 14433
rect 5632 14424 5684 14476
rect 3516 14220 3568 14272
rect 4620 14220 4672 14272
rect 5448 14288 5500 14340
rect 6736 14467 6788 14476
rect 6736 14433 6745 14467
rect 6745 14433 6779 14467
rect 6779 14433 6788 14467
rect 6736 14424 6788 14433
rect 6828 14424 6880 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7840 14560 7892 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 9036 14560 9088 14612
rect 9496 14603 9548 14612
rect 9496 14569 9505 14603
rect 9505 14569 9539 14603
rect 9539 14569 9548 14603
rect 9496 14560 9548 14569
rect 13912 14560 13964 14612
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 9312 14467 9364 14476
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 12624 14492 12676 14544
rect 16948 14560 17000 14612
rect 9312 14424 9364 14433
rect 11152 14424 11204 14476
rect 13452 14424 13504 14476
rect 13544 14467 13596 14476
rect 13544 14433 13553 14467
rect 13553 14433 13587 14467
rect 13587 14433 13596 14467
rect 13544 14424 13596 14433
rect 14924 14424 14976 14476
rect 15108 14424 15160 14476
rect 6644 14356 6696 14408
rect 8484 14356 8536 14408
rect 9588 14356 9640 14408
rect 10784 14356 10836 14408
rect 11428 14331 11480 14340
rect 11428 14297 11437 14331
rect 11437 14297 11471 14331
rect 11471 14297 11480 14331
rect 11428 14288 11480 14297
rect 12072 14356 12124 14408
rect 14372 14356 14424 14408
rect 14740 14288 14792 14340
rect 6644 14263 6696 14272
rect 6644 14229 6653 14263
rect 6653 14229 6687 14263
rect 6687 14229 6696 14263
rect 6644 14220 6696 14229
rect 11244 14220 11296 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 13452 14220 13504 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16580 14424 16632 14476
rect 16672 14424 16724 14476
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 17408 14424 17460 14476
rect 16488 14288 16540 14340
rect 17316 14220 17368 14272
rect 18144 14220 18196 14272
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 2228 14016 2280 14068
rect 5448 14059 5500 14068
rect 5448 14025 5457 14059
rect 5457 14025 5491 14059
rect 5491 14025 5500 14059
rect 5448 14016 5500 14025
rect 5632 14016 5684 14068
rect 8208 14016 8260 14068
rect 11428 14016 11480 14068
rect 15108 14059 15160 14068
rect 15108 14025 15117 14059
rect 15117 14025 15151 14059
rect 15151 14025 15160 14059
rect 15108 14016 15160 14025
rect 16580 14059 16632 14068
rect 16580 14025 16589 14059
rect 16589 14025 16623 14059
rect 16623 14025 16632 14059
rect 16580 14016 16632 14025
rect 2320 13923 2372 13932
rect 2320 13889 2329 13923
rect 2329 13889 2363 13923
rect 2363 13889 2372 13923
rect 2320 13880 2372 13889
rect 2136 13812 2188 13864
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 3424 13812 3476 13864
rect 3976 13855 4028 13864
rect 3976 13821 3985 13855
rect 3985 13821 4019 13855
rect 4019 13821 4028 13855
rect 3976 13812 4028 13821
rect 5632 13855 5684 13864
rect 5632 13821 5641 13855
rect 5641 13821 5675 13855
rect 5675 13821 5684 13855
rect 5632 13812 5684 13821
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 6644 13855 6696 13864
rect 2964 13744 3016 13796
rect 4436 13744 4488 13796
rect 6000 13787 6052 13796
rect 6000 13753 6009 13787
rect 6009 13753 6043 13787
rect 6043 13753 6052 13787
rect 6000 13744 6052 13753
rect 6644 13821 6678 13855
rect 6678 13821 6696 13855
rect 6644 13812 6696 13821
rect 11060 13812 11112 13864
rect 6736 13744 6788 13796
rect 11244 13812 11296 13864
rect 13912 13880 13964 13932
rect 17684 13948 17736 14000
rect 13452 13744 13504 13796
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 15292 13812 15344 13864
rect 15476 13855 15528 13864
rect 15476 13821 15510 13855
rect 15510 13821 15528 13855
rect 15476 13812 15528 13821
rect 16948 13812 17000 13864
rect 14740 13744 14792 13796
rect 15108 13787 15160 13796
rect 15108 13753 15117 13787
rect 15117 13753 15151 13787
rect 15151 13753 15160 13787
rect 15108 13744 15160 13753
rect 3148 13676 3200 13728
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 12624 13676 12676 13728
rect 12716 13676 12768 13728
rect 13728 13719 13780 13728
rect 13728 13685 13737 13719
rect 13737 13685 13771 13719
rect 13771 13685 13780 13719
rect 13728 13676 13780 13685
rect 14372 13676 14424 13728
rect 14924 13676 14976 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 2504 13472 2556 13524
rect 2964 13472 3016 13524
rect 4436 13515 4488 13524
rect 4436 13481 4445 13515
rect 4445 13481 4479 13515
rect 4479 13481 4488 13515
rect 4436 13472 4488 13481
rect 8944 13404 8996 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 6000 13336 6052 13388
rect 7288 13336 7340 13388
rect 8484 13379 8536 13388
rect 8484 13345 8493 13379
rect 8493 13345 8527 13379
rect 8527 13345 8536 13379
rect 8484 13336 8536 13345
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2596 13268 2648 13320
rect 3332 13268 3384 13320
rect 8208 13268 8260 13320
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 11612 13336 11664 13388
rect 10692 13268 10744 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 15108 13472 15160 13524
rect 12624 13404 12676 13456
rect 12716 13447 12768 13456
rect 12716 13413 12741 13447
rect 12741 13413 12768 13447
rect 12716 13404 12768 13413
rect 15200 13404 15252 13456
rect 13912 13379 13964 13388
rect 13912 13345 13921 13379
rect 13921 13345 13955 13379
rect 13955 13345 13964 13379
rect 13912 13336 13964 13345
rect 14004 13336 14056 13388
rect 2320 13200 2372 13252
rect 1032 13175 1084 13184
rect 1032 13141 1041 13175
rect 1041 13141 1075 13175
rect 1075 13141 1084 13175
rect 1032 13132 1084 13141
rect 6920 13132 6972 13184
rect 8668 13132 8720 13184
rect 8852 13175 8904 13184
rect 8852 13141 8861 13175
rect 8861 13141 8895 13175
rect 8895 13141 8904 13175
rect 8852 13132 8904 13141
rect 9680 13132 9732 13184
rect 10784 13200 10836 13252
rect 13544 13268 13596 13320
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 17500 13379 17552 13388
rect 17500 13345 17509 13379
rect 17509 13345 17543 13379
rect 17543 13345 17552 13379
rect 17500 13336 17552 13345
rect 18144 13515 18196 13524
rect 18144 13481 18153 13515
rect 18153 13481 18187 13515
rect 18187 13481 18196 13515
rect 18144 13472 18196 13481
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 11152 13132 11204 13184
rect 12072 13132 12124 13184
rect 12532 13132 12584 13184
rect 13728 13132 13780 13184
rect 16120 13175 16172 13184
rect 16120 13141 16129 13175
rect 16129 13141 16163 13175
rect 16163 13141 16172 13175
rect 16120 13132 16172 13141
rect 18788 13175 18840 13184
rect 18788 13141 18797 13175
rect 18797 13141 18831 13175
rect 18831 13141 18840 13175
rect 18788 13132 18840 13141
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 1860 12928 1912 12980
rect 7196 12860 7248 12912
rect 8208 12971 8260 12980
rect 8208 12937 8217 12971
rect 8217 12937 8251 12971
rect 8251 12937 8260 12971
rect 8208 12928 8260 12937
rect 8760 12928 8812 12980
rect 9220 12928 9272 12980
rect 8484 12860 8536 12912
rect 1032 12835 1084 12844
rect 1032 12801 1041 12835
rect 1041 12801 1075 12835
rect 1075 12801 1084 12835
rect 1032 12792 1084 12801
rect 3332 12835 3384 12844
rect 3332 12801 3341 12835
rect 3341 12801 3375 12835
rect 3375 12801 3384 12835
rect 3332 12792 3384 12801
rect 3056 12767 3108 12776
rect 3056 12733 3065 12767
rect 3065 12733 3099 12767
rect 3099 12733 3108 12767
rect 3056 12724 3108 12733
rect 3148 12656 3200 12708
rect 3240 12699 3292 12708
rect 3240 12665 3249 12699
rect 3249 12665 3283 12699
rect 3283 12665 3292 12699
rect 3240 12656 3292 12665
rect 3516 12767 3568 12776
rect 3516 12733 3525 12767
rect 3525 12733 3559 12767
rect 3559 12733 3568 12767
rect 3516 12724 3568 12733
rect 7104 12767 7156 12776
rect 7104 12733 7113 12767
rect 7113 12733 7147 12767
rect 7147 12733 7156 12767
rect 7104 12724 7156 12733
rect 7288 12724 7340 12776
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8484 12767 8536 12776
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 8484 12724 8536 12733
rect 10508 12928 10560 12980
rect 10692 12860 10744 12912
rect 11336 12792 11388 12844
rect 11152 12724 11204 12776
rect 11520 12724 11572 12776
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 3976 12656 4028 12708
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2596 12588 2648 12640
rect 6460 12656 6512 12708
rect 8852 12656 8904 12708
rect 12072 12860 12124 12912
rect 12164 12724 12216 12776
rect 12624 12724 12676 12776
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 12900 12835 12952 12844
rect 12900 12801 12909 12835
rect 12909 12801 12943 12835
rect 12943 12801 12952 12835
rect 12900 12792 12952 12801
rect 13084 12971 13136 12980
rect 13084 12937 13093 12971
rect 13093 12937 13127 12971
rect 13127 12937 13136 12971
rect 13084 12928 13136 12937
rect 14004 12971 14056 12980
rect 14004 12937 14013 12971
rect 14013 12937 14047 12971
rect 14047 12937 14056 12971
rect 14004 12928 14056 12937
rect 18420 12971 18472 12980
rect 18420 12937 18429 12971
rect 18429 12937 18463 12971
rect 18463 12937 18472 12971
rect 18420 12928 18472 12937
rect 18604 12928 18656 12980
rect 16672 12860 16724 12912
rect 14188 12792 14240 12844
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 14924 12792 14976 12844
rect 15292 12792 15344 12844
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 13820 12767 13872 12776
rect 13820 12733 13829 12767
rect 13829 12733 13863 12767
rect 13863 12733 13872 12767
rect 13820 12724 13872 12733
rect 9680 12588 9732 12640
rect 11428 12588 11480 12640
rect 12440 12631 12492 12640
rect 12440 12597 12449 12631
rect 12449 12597 12483 12631
rect 12483 12597 12492 12631
rect 12440 12588 12492 12597
rect 12532 12588 12584 12640
rect 14372 12767 14424 12776
rect 14372 12733 14381 12767
rect 14381 12733 14415 12767
rect 14415 12733 14424 12767
rect 14372 12724 14424 12733
rect 15108 12656 15160 12708
rect 16488 12656 16540 12708
rect 18788 12724 18840 12776
rect 16856 12588 16908 12640
rect 17500 12588 17552 12640
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 1860 12384 1912 12436
rect 1584 12316 1636 12368
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 6828 12427 6880 12436
rect 6828 12393 6837 12427
rect 6837 12393 6871 12427
rect 6871 12393 6880 12427
rect 6828 12384 6880 12393
rect 1676 12248 1728 12300
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 3056 12180 3108 12232
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4712 12359 4764 12368
rect 4712 12325 4721 12359
rect 4721 12325 4755 12359
rect 4755 12325 4764 12359
rect 4712 12316 4764 12325
rect 4988 12248 5040 12300
rect 6000 12316 6052 12368
rect 6920 12359 6972 12368
rect 6920 12325 6929 12359
rect 6929 12325 6963 12359
rect 6963 12325 6972 12359
rect 6920 12316 6972 12325
rect 7380 12359 7432 12368
rect 7380 12325 7389 12359
rect 7389 12325 7423 12359
rect 7423 12325 7432 12359
rect 7380 12316 7432 12325
rect 5540 12291 5592 12300
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 5816 12248 5868 12300
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 7104 12248 7156 12300
rect 7288 12291 7340 12300
rect 7288 12257 7297 12291
rect 7297 12257 7331 12291
rect 7331 12257 7340 12291
rect 7288 12248 7340 12257
rect 8484 12316 8536 12368
rect 9496 12384 9548 12436
rect 8668 12291 8720 12300
rect 8668 12257 8686 12291
rect 8686 12257 8720 12291
rect 8668 12248 8720 12257
rect 9128 12248 9180 12300
rect 9680 12316 9732 12368
rect 11244 12316 11296 12368
rect 13912 12359 13964 12368
rect 13912 12325 13921 12359
rect 13921 12325 13955 12359
rect 13955 12325 13964 12359
rect 13912 12316 13964 12325
rect 9772 12248 9824 12300
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 3148 12044 3200 12096
rect 4528 12044 4580 12096
rect 11428 12291 11480 12300
rect 11428 12257 11437 12291
rect 11437 12257 11471 12291
rect 11471 12257 11480 12291
rect 11428 12248 11480 12257
rect 11520 12248 11572 12300
rect 13636 12248 13688 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 17500 12291 17552 12300
rect 17500 12257 17509 12291
rect 17509 12257 17543 12291
rect 17543 12257 17552 12291
rect 17500 12248 17552 12257
rect 12072 12180 12124 12232
rect 12532 12112 12584 12164
rect 5816 12044 5868 12096
rect 7288 12044 7340 12096
rect 7656 12044 7708 12096
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 11428 12087 11480 12096
rect 11428 12053 11437 12087
rect 11437 12053 11471 12087
rect 11471 12053 11480 12087
rect 11428 12044 11480 12053
rect 15016 12044 15068 12096
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 3148 11840 3200 11892
rect 3424 11840 3476 11892
rect 4068 11840 4120 11892
rect 4252 11840 4304 11892
rect 5540 11840 5592 11892
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 9680 11840 9732 11892
rect 12532 11840 12584 11892
rect 2320 11772 2372 11824
rect 3240 11747 3292 11756
rect 3240 11713 3249 11747
rect 3249 11713 3283 11747
rect 3283 11713 3292 11747
rect 3240 11704 3292 11713
rect 3976 11815 4028 11824
rect 3976 11781 3985 11815
rect 3985 11781 4019 11815
rect 4019 11781 4028 11815
rect 3976 11772 4028 11781
rect 4712 11772 4764 11824
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 6460 11747 6512 11756
rect 6460 11713 6469 11747
rect 6469 11713 6503 11747
rect 6503 11713 6512 11747
rect 6460 11704 6512 11713
rect 4068 11568 4120 11620
rect 6000 11568 6052 11620
rect 7288 11636 7340 11688
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 10968 11636 11020 11688
rect 11428 11636 11480 11688
rect 12808 11704 12860 11756
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 13820 11840 13872 11892
rect 15936 11840 15988 11892
rect 13268 11772 13320 11824
rect 13452 11704 13504 11756
rect 13636 11636 13688 11688
rect 16396 11704 16448 11756
rect 10600 11500 10652 11552
rect 12072 11500 12124 11552
rect 12992 11500 13044 11552
rect 14924 11636 14976 11688
rect 15200 11636 15252 11688
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 14188 11500 14240 11552
rect 15016 11500 15068 11552
rect 15292 11500 15344 11552
rect 15936 11543 15988 11552
rect 15936 11509 15945 11543
rect 15945 11509 15979 11543
rect 15979 11509 15988 11543
rect 15936 11500 15988 11509
rect 16488 11500 16540 11552
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 2228 11296 2280 11348
rect 3240 11296 3292 11348
rect 4988 11296 5040 11348
rect 6000 11339 6052 11348
rect 6000 11305 6009 11339
rect 6009 11305 6043 11339
rect 6043 11305 6052 11339
rect 6000 11296 6052 11305
rect 3976 11160 4028 11212
rect 8576 11228 8628 11280
rect 4528 11203 4580 11212
rect 4528 11169 4562 11203
rect 4562 11169 4580 11203
rect 4528 11160 4580 11169
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 10416 11228 10468 11280
rect 13084 11228 13136 11280
rect 17408 11228 17460 11280
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 9404 11203 9456 11212
rect 9404 11169 9413 11203
rect 9413 11169 9447 11203
rect 9447 11169 9456 11203
rect 9404 11160 9456 11169
rect 9588 11203 9640 11212
rect 9588 11169 9597 11203
rect 9597 11169 9631 11203
rect 9631 11169 9640 11203
rect 9588 11160 9640 11169
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 13268 11203 13320 11212
rect 13268 11169 13277 11203
rect 13277 11169 13311 11203
rect 13311 11169 13320 11203
rect 13268 11160 13320 11169
rect 15108 11160 15160 11212
rect 16396 11160 16448 11212
rect 17868 11228 17920 11280
rect 14188 11092 14240 11144
rect 8944 11024 8996 11076
rect 9312 11024 9364 11076
rect 10232 11024 10284 11076
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 16672 11092 16724 11101
rect 17224 11024 17276 11076
rect 17408 10956 17460 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 13084 10752 13136 10804
rect 14924 10752 14976 10804
rect 10968 10684 11020 10736
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 16488 10684 16540 10736
rect 7932 10548 7984 10600
rect 9588 10548 9640 10600
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 10784 10591 10836 10600
rect 10784 10557 10793 10591
rect 10793 10557 10827 10591
rect 10827 10557 10836 10591
rect 10784 10548 10836 10557
rect 12716 10591 12768 10600
rect 12716 10557 12725 10591
rect 12725 10557 12759 10591
rect 12759 10557 12768 10591
rect 12716 10548 12768 10557
rect 13268 10548 13320 10600
rect 14096 10591 14148 10600
rect 14096 10557 14105 10591
rect 14105 10557 14139 10591
rect 14139 10557 14148 10591
rect 14096 10548 14148 10557
rect 14372 10616 14424 10668
rect 15016 10616 15068 10668
rect 9680 10412 9732 10464
rect 13268 10412 13320 10464
rect 13360 10455 13412 10464
rect 13360 10421 13369 10455
rect 13369 10421 13403 10455
rect 13403 10421 13412 10455
rect 13360 10412 13412 10421
rect 14004 10480 14056 10532
rect 15200 10548 15252 10600
rect 16396 10591 16448 10600
rect 16396 10557 16405 10591
rect 16405 10557 16439 10591
rect 16439 10557 16448 10591
rect 16396 10548 16448 10557
rect 16580 10591 16632 10600
rect 16580 10557 16589 10591
rect 16589 10557 16623 10591
rect 16623 10557 16632 10591
rect 16580 10548 16632 10557
rect 15108 10480 15160 10532
rect 17224 10548 17276 10600
rect 18052 10523 18104 10532
rect 18052 10489 18061 10523
rect 18061 10489 18095 10523
rect 18095 10489 18104 10523
rect 18052 10480 18104 10489
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 11152 10208 11204 10260
rect 9588 10140 9640 10192
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 10784 10140 10836 10192
rect 10416 10115 10468 10124
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 10876 10072 10928 10124
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 13452 10208 13504 10260
rect 13360 10140 13412 10192
rect 10692 10004 10744 10056
rect 10048 9979 10100 9988
rect 10048 9945 10057 9979
rect 10057 9945 10091 9979
rect 10091 9945 10100 9979
rect 10048 9936 10100 9945
rect 10140 9868 10192 9920
rect 11336 9936 11388 9988
rect 12992 9936 13044 9988
rect 14096 10072 14148 10124
rect 18052 10208 18104 10260
rect 15200 10183 15252 10192
rect 15200 10149 15209 10183
rect 15209 10149 15243 10183
rect 15243 10149 15252 10183
rect 15200 10140 15252 10149
rect 13912 10004 13964 10056
rect 14924 10072 14976 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 16120 10072 16172 10124
rect 16580 10004 16632 10056
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 17868 10004 17920 10056
rect 10784 9911 10836 9920
rect 10784 9877 10793 9911
rect 10793 9877 10827 9911
rect 10827 9877 10836 9911
rect 10784 9868 10836 9877
rect 11612 9911 11664 9920
rect 11612 9877 11621 9911
rect 11621 9877 11655 9911
rect 11655 9877 11664 9911
rect 11612 9868 11664 9877
rect 13912 9911 13964 9920
rect 13912 9877 13921 9911
rect 13921 9877 13955 9911
rect 13955 9877 13964 9911
rect 13912 9868 13964 9877
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 15292 9936 15344 9988
rect 16120 9868 16172 9920
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 9680 9664 9732 9716
rect 10692 9664 10744 9716
rect 13176 9664 13228 9716
rect 15292 9664 15344 9716
rect 8852 9639 8904 9648
rect 8852 9605 8861 9639
rect 8861 9605 8895 9639
rect 8895 9605 8904 9639
rect 8852 9596 8904 9605
rect 9496 9596 9548 9648
rect 9772 9596 9824 9648
rect 9956 9528 10008 9580
rect 10324 9528 10376 9580
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 10784 9460 10836 9512
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 12532 9528 12584 9580
rect 12992 9528 13044 9580
rect 10876 9460 10928 9469
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 10048 9392 10100 9444
rect 10600 9435 10652 9444
rect 10600 9401 10609 9435
rect 10609 9401 10643 9435
rect 10643 9401 10652 9435
rect 10600 9392 10652 9401
rect 12256 9503 12308 9512
rect 12256 9469 12265 9503
rect 12265 9469 12299 9503
rect 12299 9469 12308 9503
rect 12256 9460 12308 9469
rect 12900 9460 12952 9512
rect 13268 9528 13320 9580
rect 13820 9596 13872 9648
rect 14280 9596 14332 9648
rect 15200 9596 15252 9648
rect 15844 9596 15896 9648
rect 16028 9596 16080 9648
rect 16948 9596 17000 9648
rect 14096 9528 14148 9580
rect 14188 9528 14240 9580
rect 15752 9528 15804 9580
rect 17684 9528 17736 9580
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 13636 9460 13688 9512
rect 13728 9392 13780 9444
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10324 9324 10376 9376
rect 10508 9324 10560 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 12624 9324 12676 9376
rect 13084 9324 13136 9376
rect 13636 9324 13688 9376
rect 15016 9460 15068 9512
rect 15844 9503 15896 9512
rect 15844 9469 15853 9503
rect 15853 9469 15887 9503
rect 15887 9469 15896 9503
rect 15844 9460 15896 9469
rect 16580 9460 16632 9512
rect 14464 9392 14516 9444
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 15016 9324 15068 9376
rect 16120 9324 16172 9376
rect 16488 9324 16540 9376
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 10416 9120 10468 9172
rect 9404 9052 9456 9104
rect 11336 9120 11388 9172
rect 12900 9163 12952 9172
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 13636 9163 13688 9172
rect 13636 9129 13645 9163
rect 13645 9129 13679 9163
rect 13679 9129 13688 9163
rect 13636 9120 13688 9129
rect 13728 9120 13780 9172
rect 11244 9052 11296 9104
rect 14464 9052 14516 9104
rect 9220 9027 9272 9036
rect 9220 8993 9229 9027
rect 9229 8993 9263 9027
rect 9263 8993 9272 9027
rect 9220 8984 9272 8993
rect 10324 8984 10376 9036
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 14188 8984 14240 9036
rect 14372 8984 14424 9036
rect 13268 8959 13320 8968
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 13544 8916 13596 8968
rect 13728 8916 13780 8968
rect 14004 8959 14056 8968
rect 14004 8925 14013 8959
rect 14013 8925 14047 8959
rect 14047 8925 14056 8959
rect 14004 8916 14056 8925
rect 14464 8916 14516 8968
rect 14740 9027 14792 9036
rect 14740 8993 14749 9027
rect 14749 8993 14783 9027
rect 14783 8993 14792 9027
rect 14740 8984 14792 8993
rect 15384 8984 15436 9036
rect 16028 9120 16080 9172
rect 16212 9120 16264 9172
rect 16580 9163 16632 9172
rect 16580 9129 16589 9163
rect 16589 9129 16623 9163
rect 16623 9129 16632 9163
rect 16580 9120 16632 9129
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 17684 9120 17736 9172
rect 18236 9120 18288 9172
rect 15292 8916 15344 8968
rect 16028 8984 16080 9036
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 17408 8984 17460 9036
rect 17684 9027 17736 9036
rect 17684 8993 17693 9027
rect 17693 8993 17727 9027
rect 17727 8993 17736 9027
rect 17684 8984 17736 8993
rect 17776 8984 17828 9036
rect 18052 9052 18104 9104
rect 17960 9027 18012 9036
rect 17960 8993 17969 9027
rect 17969 8993 18003 9027
rect 18003 8993 18012 9027
rect 17960 8984 18012 8993
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 18420 9027 18472 9036
rect 18420 8993 18429 9027
rect 18429 8993 18463 9027
rect 18463 8993 18472 9027
rect 18420 8984 18472 8993
rect 16120 8916 16172 8968
rect 16672 8959 16724 8968
rect 16672 8925 16681 8959
rect 16681 8925 16715 8959
rect 16715 8925 16724 8959
rect 16672 8916 16724 8925
rect 9864 8848 9916 8900
rect 12440 8848 12492 8900
rect 13084 8848 13136 8900
rect 7932 8823 7984 8832
rect 7932 8789 7941 8823
rect 7941 8789 7975 8823
rect 7975 8789 7984 8823
rect 7932 8780 7984 8789
rect 11796 8780 11848 8832
rect 16212 8848 16264 8900
rect 15292 8780 15344 8832
rect 16028 8780 16080 8832
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 16304 8780 16356 8832
rect 17960 8848 18012 8900
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 13176 8576 13228 8628
rect 13820 8576 13872 8628
rect 15936 8576 15988 8628
rect 16304 8576 16356 8628
rect 16488 8576 16540 8628
rect 8576 8508 8628 8560
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 11704 8440 11756 8492
rect 8852 8372 8904 8424
rect 14188 8508 14240 8560
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 12164 8415 12216 8424
rect 12164 8381 12173 8415
rect 12173 8381 12207 8415
rect 12207 8381 12216 8415
rect 12164 8372 12216 8381
rect 12440 8372 12492 8424
rect 10784 8304 10836 8356
rect 13636 8372 13688 8424
rect 14096 8372 14148 8424
rect 14740 8440 14792 8492
rect 13084 8347 13136 8356
rect 13084 8313 13093 8347
rect 13093 8313 13127 8347
rect 13127 8313 13136 8347
rect 13084 8304 13136 8313
rect 13728 8347 13780 8356
rect 13728 8313 13737 8347
rect 13737 8313 13771 8347
rect 13771 8313 13780 8347
rect 13728 8304 13780 8313
rect 13912 8347 13964 8356
rect 13912 8313 13921 8347
rect 13921 8313 13955 8347
rect 13955 8313 13964 8347
rect 13912 8304 13964 8313
rect 14464 8372 14516 8424
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 17040 8508 17092 8560
rect 17500 8508 17552 8560
rect 17868 8508 17920 8560
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 15200 8415 15252 8424
rect 15200 8381 15209 8415
rect 15209 8381 15243 8415
rect 15243 8381 15252 8415
rect 15200 8372 15252 8381
rect 15292 8415 15344 8424
rect 15292 8381 15301 8415
rect 15301 8381 15335 8415
rect 15335 8381 15344 8415
rect 15292 8372 15344 8381
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 15568 8415 15620 8424
rect 15568 8381 15577 8415
rect 15577 8381 15611 8415
rect 15611 8381 15620 8415
rect 15568 8372 15620 8381
rect 15660 8415 15712 8424
rect 15660 8381 15669 8415
rect 15669 8381 15703 8415
rect 15703 8381 15712 8415
rect 15660 8372 15712 8381
rect 15476 8304 15528 8356
rect 16120 8372 16172 8424
rect 17776 8440 17828 8492
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 17408 8372 17460 8424
rect 17316 8304 17368 8356
rect 18420 8372 18472 8424
rect 11980 8279 12032 8288
rect 11980 8245 11989 8279
rect 11989 8245 12023 8279
rect 12023 8245 12032 8279
rect 11980 8236 12032 8245
rect 13268 8236 13320 8288
rect 17500 8236 17552 8288
rect 17592 8279 17644 8288
rect 17592 8245 17601 8279
rect 17601 8245 17635 8279
rect 17635 8245 17644 8279
rect 17592 8236 17644 8245
rect 18236 8236 18288 8288
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 10232 8032 10284 8084
rect 10600 8032 10652 8084
rect 12164 8075 12216 8084
rect 12164 8041 12173 8075
rect 12173 8041 12207 8075
rect 12207 8041 12216 8075
rect 12164 8032 12216 8041
rect 12440 8032 12492 8084
rect 9588 7964 9640 8016
rect 10324 7964 10376 8016
rect 10968 7964 11020 8016
rect 11980 7828 12032 7880
rect 12532 7939 12584 7948
rect 12532 7905 12541 7939
rect 12541 7905 12575 7939
rect 12575 7905 12584 7939
rect 12532 7896 12584 7905
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 12808 7896 12860 7905
rect 13360 8032 13412 8084
rect 14924 8032 14976 8084
rect 15660 8032 15712 8084
rect 13452 7896 13504 7948
rect 15200 7964 15252 8016
rect 14464 7939 14516 7948
rect 14464 7905 14473 7939
rect 14473 7905 14507 7939
rect 14507 7905 14516 7939
rect 14464 7896 14516 7905
rect 13636 7828 13688 7880
rect 14924 7896 14976 7948
rect 17040 7939 17092 7948
rect 17040 7905 17049 7939
rect 17049 7905 17083 7939
rect 17083 7905 17092 7939
rect 17040 7896 17092 7905
rect 15016 7828 15068 7880
rect 15292 7828 15344 7880
rect 15936 7828 15988 7880
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 17500 7896 17552 7948
rect 17592 7896 17644 7948
rect 17960 7939 18012 7948
rect 17960 7905 17969 7939
rect 17969 7905 18003 7939
rect 18003 7905 18012 7939
rect 17960 7896 18012 7905
rect 10232 7692 10284 7744
rect 13268 7692 13320 7744
rect 13728 7692 13780 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 17500 7692 17552 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 9680 7352 9732 7404
rect 10600 7352 10652 7404
rect 12808 7488 12860 7540
rect 14280 7488 14332 7540
rect 17224 7488 17276 7540
rect 18052 7488 18104 7540
rect 13820 7352 13872 7404
rect 15936 7420 15988 7472
rect 9036 7284 9088 7336
rect 10968 7327 11020 7336
rect 10968 7293 10977 7327
rect 10977 7293 11011 7327
rect 11011 7293 11020 7327
rect 10968 7284 11020 7293
rect 11704 7284 11756 7336
rect 8392 7259 8444 7268
rect 8392 7225 8401 7259
rect 8401 7225 8435 7259
rect 8435 7225 8444 7259
rect 8392 7216 8444 7225
rect 10508 7148 10560 7200
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 13084 7216 13136 7268
rect 14004 7284 14056 7336
rect 14464 7327 14516 7336
rect 14464 7293 14473 7327
rect 14473 7293 14507 7327
rect 14507 7293 14516 7327
rect 15752 7352 15804 7404
rect 14464 7284 14516 7293
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 15844 7284 15896 7336
rect 17500 7395 17552 7404
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 16580 7284 16632 7336
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 13176 7148 13228 7200
rect 14004 7148 14056 7200
rect 15108 7216 15160 7268
rect 15292 7216 15344 7268
rect 14280 7148 14332 7200
rect 15476 7148 15528 7200
rect 15568 7148 15620 7200
rect 15844 7191 15896 7200
rect 15844 7157 15853 7191
rect 15853 7157 15887 7191
rect 15887 7157 15896 7191
rect 15844 7148 15896 7157
rect 16856 7148 16908 7200
rect 17408 7148 17460 7200
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 10140 6944 10192 6996
rect 10600 6944 10652 6996
rect 13176 6944 13228 6996
rect 13544 6944 13596 6996
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 9404 6851 9456 6860
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 9956 6919 10008 6928
rect 9956 6885 9965 6919
rect 9965 6885 9999 6919
rect 9999 6885 10008 6919
rect 9956 6876 10008 6885
rect 10968 6876 11020 6928
rect 13452 6876 13504 6928
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 9588 6808 9640 6860
rect 9036 6672 9088 6724
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 10692 6808 10744 6860
rect 10784 6851 10836 6860
rect 10784 6817 10793 6851
rect 10793 6817 10827 6851
rect 10827 6817 10836 6851
rect 10784 6808 10836 6817
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 12624 6808 12676 6860
rect 12716 6808 12768 6860
rect 11152 6740 11204 6792
rect 10692 6672 10744 6724
rect 11244 6672 11296 6724
rect 12532 6672 12584 6724
rect 12716 6672 12768 6724
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14372 6851 14424 6860
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 15384 6876 15436 6928
rect 15292 6808 15344 6860
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 16028 6944 16080 6996
rect 16672 6919 16724 6928
rect 16672 6885 16681 6919
rect 16681 6885 16715 6919
rect 16715 6885 16724 6919
rect 16672 6876 16724 6885
rect 15016 6740 15068 6792
rect 15200 6740 15252 6792
rect 9496 6604 9548 6656
rect 10968 6647 11020 6656
rect 10968 6613 10977 6647
rect 10977 6613 11011 6647
rect 11011 6613 11020 6647
rect 10968 6604 11020 6613
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 13728 6604 13780 6656
rect 14464 6647 14516 6656
rect 14464 6613 14473 6647
rect 14473 6613 14507 6647
rect 14507 6613 14516 6647
rect 14464 6604 14516 6613
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 17316 6604 17368 6656
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 9404 6400 9456 6452
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 14648 6400 14700 6452
rect 11060 6375 11112 6384
rect 11060 6341 11069 6375
rect 11069 6341 11103 6375
rect 11103 6341 11112 6375
rect 11060 6332 11112 6341
rect 11152 6332 11204 6384
rect 14464 6332 14516 6384
rect 15200 6332 15252 6384
rect 10692 6264 10744 6316
rect 9956 6196 10008 6248
rect 10968 6196 11020 6248
rect 12532 6264 12584 6316
rect 15844 6400 15896 6452
rect 17316 6400 17368 6452
rect 15476 6332 15528 6384
rect 13544 6196 13596 6248
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 14188 6239 14240 6248
rect 14188 6205 14197 6239
rect 14197 6205 14231 6239
rect 14231 6205 14240 6239
rect 14188 6196 14240 6205
rect 15660 6264 15712 6316
rect 15752 6264 15804 6316
rect 14924 6196 14976 6248
rect 15108 6196 15160 6248
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 16580 6196 16632 6248
rect 16764 6128 16816 6180
rect 16948 6196 17000 6248
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 17316 6196 17368 6248
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 9680 5788 9732 5840
rect 9496 5720 9548 5772
rect 11060 5788 11112 5840
rect 10968 5720 11020 5772
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 13636 5516 13688 5568
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 9680 5312 9732 5364
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 10232 5108 10284 5160
rect 11244 5083 11296 5092
rect 11244 5049 11278 5083
rect 11278 5049 11296 5083
rect 11244 5040 11296 5049
rect 11612 5040 11664 5092
rect 11060 4972 11112 5024
rect 16120 4972 16172 5024
rect 18604 4972 18656 5024
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 3700 4088 3752 4140
rect 7932 4088 7984 4140
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 6184 3680 6236 3732
rect 8668 3680 8720 3732
rect 1216 3612 1268 3664
rect 8392 3612 8444 3664
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 846 19600 902 20000
rect 2502 19600 2558 20000
rect 4158 19600 4214 20000
rect 5814 19600 5870 20000
rect 7470 19600 7526 20000
rect 9126 19600 9182 20000
rect 10782 19600 10838 20000
rect 10888 19638 11100 19666
rect 860 18834 888 19600
rect 2516 18834 2544 19600
rect 4172 18834 4200 19600
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 5828 18834 5856 19600
rect 7484 18834 7512 19600
rect 9140 18834 9168 19600
rect 10796 19530 10824 19600
rect 10888 19530 10916 19638
rect 10796 19502 10916 19530
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 848 18828 900 18834
rect 848 18770 900 18776
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 9128 18828 9180 18834
rect 9128 18770 9180 18776
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 2755 18459 3063 18468
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4172 17746 4200 18158
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 1872 16046 1900 17070
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16726 2452 16934
rect 3712 16726 3740 17070
rect 2412 16720 2464 16726
rect 2412 16662 2464 16668
rect 3700 16720 3752 16726
rect 3700 16662 3752 16668
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15638 1716 15846
rect 1676 15632 1728 15638
rect 1676 15574 1728 15580
rect 2056 15552 2084 16526
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3516 16448 3568 16454
rect 3516 16390 3568 16396
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 3528 16182 3556 16390
rect 3516 16176 3568 16182
rect 3516 16118 3568 16124
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 2136 15564 2188 15570
rect 2056 15524 2136 15552
rect 1676 15088 1728 15094
rect 1676 15030 1728 15036
rect 1688 13394 1716 15030
rect 2056 14482 2084 15524
rect 2136 15506 2188 15512
rect 2332 15162 2360 15846
rect 2608 15570 2636 15846
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2792 15502 2820 15982
rect 2884 15502 2912 16050
rect 3528 16046 3556 16118
rect 3620 16046 3648 16458
rect 3896 16454 3924 17070
rect 4172 16794 4200 17682
rect 4356 17338 4384 17682
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4172 16658 4200 16730
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3988 16250 4016 16594
rect 4264 16538 4292 17138
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4172 16522 4292 16538
rect 4160 16516 4292 16522
rect 4212 16510 4292 16516
rect 4160 16458 4212 16464
rect 3976 16244 4028 16250
rect 3976 16186 4028 16192
rect 3516 16040 3568 16046
rect 3516 15982 3568 15988
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15502 3004 15914
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 15570 3372 15846
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2332 15026 2360 15098
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2136 14816 2188 14822
rect 2136 14758 2188 14764
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2148 13870 2176 14758
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2240 14074 2268 14418
rect 2228 14068 2280 14074
rect 2228 14010 2280 14016
rect 2332 13938 2360 14962
rect 2424 14890 2452 15302
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 3160 15162 3188 15438
rect 3240 15428 3292 15434
rect 3240 15370 3292 15376
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3252 14890 3280 15370
rect 2412 14884 2464 14890
rect 2412 14826 2464 14832
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3344 14822 3372 15506
rect 4172 15502 4200 16458
rect 4448 15706 4476 16594
rect 4632 16182 4660 17070
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 5460 16250 5488 17546
rect 5736 17202 5764 18022
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5828 17134 5856 17478
rect 6288 17134 6316 18022
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4632 15570 4660 16118
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3528 14278 3556 15098
rect 4172 15026 4200 15438
rect 5460 15366 5488 16050
rect 5736 16046 5764 16526
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 5724 16040 5776 16046
rect 5724 15982 5776 15988
rect 5828 15502 5856 16390
rect 6472 16046 6500 17614
rect 6932 17610 6960 18566
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 7024 17270 7052 18362
rect 7208 18170 7236 18702
rect 8024 18692 8076 18698
rect 8024 18634 8076 18640
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 7288 18216 7340 18222
rect 7208 18164 7288 18170
rect 7208 18158 7340 18164
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7208 18142 7328 18158
rect 7472 18148 7524 18154
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7116 17338 7144 18022
rect 7208 17746 7236 18142
rect 7472 18090 7524 18096
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7380 18080 7432 18086
rect 7380 18022 7432 18028
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7024 16454 7052 17206
rect 7208 16998 7236 17478
rect 7300 17202 7328 18022
rect 7392 17882 7420 18022
rect 7484 17882 7512 18090
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7576 17678 7604 18158
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17746 7788 18022
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7484 17542 7512 17614
rect 7760 17610 7788 17682
rect 7748 17604 7800 17610
rect 7748 17546 7800 17552
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 7024 16232 7052 16390
rect 6932 16204 7052 16232
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 4080 14482 4476 14498
rect 4068 14476 4488 14482
rect 4120 14470 4436 14476
rect 4068 14418 4120 14424
rect 4436 14418 4488 14424
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1032 13184 1084 13190
rect 1032 13126 1084 13132
rect 1044 12850 1072 13126
rect 1032 12844 1084 12850
rect 1032 12786 1084 12792
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12374 1624 12582
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1688 12306 1716 13330
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 2332 13258 2360 13874
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 2516 13530 2544 13806
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2976 13530 3004 13738
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1872 12442 1900 12922
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2240 11354 2268 12174
rect 2332 11830 2360 13194
rect 2608 12646 2636 13262
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 3056 12776 3108 12782
rect 3056 12718 3108 12724
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12102 2636 12582
rect 3068 12238 3096 12718
rect 3160 12714 3188 13670
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3344 12850 3372 13262
rect 3332 12844 3384 12850
rect 3332 12786 3384 12792
rect 3148 12708 3200 12714
rect 3148 12650 3200 12656
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 3160 11898 3188 12038
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 3252 11762 3280 12650
rect 3436 11898 3464 13806
rect 3528 12782 3556 14214
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3516 12776 3568 12782
rect 3516 12718 3568 12724
rect 3988 12714 4016 13806
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 4080 12442 4108 14418
rect 5460 14346 5488 15302
rect 6184 15156 6236 15162
rect 6184 15098 6236 15104
rect 6196 14890 6224 15098
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6196 14550 6224 14826
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4448 13530 4476 13738
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4632 13394 4660 14214
rect 5460 14074 5488 14282
rect 5644 14074 5672 14418
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5644 13870 5672 14010
rect 6380 13938 6408 14894
rect 6656 14414 6684 15914
rect 6932 15706 6960 16204
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6748 14482 6776 15506
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6644 14408 6696 14414
rect 6644 14350 6696 14356
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6656 13870 6684 14214
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6748 13802 6776 14418
rect 6000 13796 6052 13802
rect 6000 13738 6052 13744
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4264 11898 4292 12242
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 3424 11892 3476 11898
rect 3424 11834 3476 11840
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3252 11354 3280 11698
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3988 11218 4016 11766
rect 4080 11626 4108 11834
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4540 11218 4568 12038
rect 4724 11830 4752 12310
rect 5828 12306 5856 13670
rect 6012 13394 6040 13738
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6012 12374 6040 13330
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 5000 11762 5028 12242
rect 5552 11898 5580 12242
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11354 5028 11698
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5828 11218 5856 12038
rect 6472 11762 6500 12650
rect 6840 12442 6868 14418
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6932 12374 6960 13126
rect 7024 12434 7052 16050
rect 7116 15570 7144 16050
rect 7208 15910 7236 16934
rect 7392 16726 7420 17070
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7852 15994 7880 17478
rect 7944 17338 7972 17478
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7944 16182 7972 17274
rect 8036 16726 8064 18634
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 8680 17746 8708 18566
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8864 17882 8892 18090
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8024 16720 8076 16726
rect 8024 16662 8076 16668
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 8116 16040 8168 16046
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7104 14884 7156 14890
rect 7104 14826 7156 14832
rect 7116 12782 7144 14826
rect 7208 14482 7236 15846
rect 7392 15706 7420 15982
rect 7852 15966 7972 15994
rect 8116 15982 8168 15988
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7288 15632 7340 15638
rect 7288 15574 7340 15580
rect 7300 15366 7328 15574
rect 7484 15450 7512 15642
rect 7392 15422 7512 15450
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7116 12617 7144 12718
rect 7102 12608 7158 12617
rect 7208 12594 7236 12854
rect 7300 12782 7328 13330
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7208 12566 7328 12594
rect 7102 12543 7158 12552
rect 7024 12406 7144 12434
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 7116 12306 7144 12406
rect 7300 12306 7328 12566
rect 7392 12374 7420 15422
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7852 14618 7880 15438
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7024 11898 7052 12242
rect 7668 12102 7696 12718
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 7300 11694 7328 12038
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6012 11354 6040 11562
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 7944 10606 7972 15966
rect 8128 15450 8156 15982
rect 8220 15570 8248 16390
rect 8404 15978 8432 17478
rect 8588 17270 8616 17682
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8680 17066 8708 17682
rect 8956 17610 8984 17682
rect 9140 17678 9168 18158
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8956 17338 8984 17546
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8404 15570 8432 15914
rect 8956 15570 8984 17274
rect 9140 16046 9168 17614
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 17202 9352 17478
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8312 15450 8340 15506
rect 8128 15422 8340 15450
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 8036 14618 8064 15302
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8220 14074 8248 15422
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8496 13394 8524 14350
rect 8956 13462 8984 15506
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 9048 14618 9076 15302
rect 9140 14958 9168 15982
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9232 15706 9260 15914
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 9416 15570 9444 18566
rect 10244 18222 10272 18566
rect 10416 18352 10468 18358
rect 10416 18294 10468 18300
rect 9680 18216 9732 18222
rect 9508 18164 9680 18170
rect 9508 18158 9732 18164
rect 10232 18216 10284 18222
rect 10284 18164 10364 18170
rect 10232 18158 10364 18164
rect 9508 18142 9720 18158
rect 10244 18142 10364 18158
rect 9508 17746 9536 18142
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9508 16658 9536 17682
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 8944 13456 8996 13462
rect 8772 13416 8944 13444
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8220 12986 8248 13262
rect 8208 12980 8260 12986
rect 8208 12922 8260 12928
rect 8496 12918 8524 13330
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8496 12374 8524 12718
rect 8484 12368 8536 12374
rect 8484 12310 8536 12316
rect 8588 11286 8616 13330
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8680 12306 8708 13126
rect 8772 12986 8800 13416
rect 8944 13398 8996 13404
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8864 12714 8892 13126
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 9140 12306 9168 13262
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9232 12102 9260 12922
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 9324 11218 9352 14418
rect 9416 11218 9444 15506
rect 9508 15434 9536 16594
rect 9600 15570 9628 17138
rect 9692 17134 9720 18022
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 17134 10180 17682
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9692 15706 9720 16730
rect 10048 16652 10100 16658
rect 10048 16594 10100 16600
rect 10060 16250 10088 16594
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9496 14884 9548 14890
rect 9496 14826 9548 14832
rect 9508 14618 9536 14826
rect 9496 14612 9548 14618
rect 9496 14554 9548 14560
rect 9600 14414 9628 15506
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12442 9536 13262
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12730 9720 13126
rect 9600 12702 9720 12730
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9600 11370 9628 12702
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12434 9720 12582
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 10244 12434 10272 18022
rect 10336 17202 10364 18142
rect 10428 17814 10456 18294
rect 10520 18222 10548 18906
rect 11072 18834 11100 19638
rect 12438 19600 12494 20000
rect 14094 19600 14150 20000
rect 15750 19600 15806 20000
rect 17406 19600 17462 20000
rect 19062 19600 19118 20000
rect 12452 18834 12480 19600
rect 14108 18834 14136 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 15764 18834 15792 19600
rect 17420 18834 17448 19600
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10428 17270 10456 17750
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10416 17128 10468 17134
rect 10520 17116 10548 18158
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 10468 17088 10548 17116
rect 10416 17070 10468 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10336 16697 10364 16934
rect 10322 16688 10378 16697
rect 10322 16623 10378 16632
rect 9692 12406 9812 12434
rect 10244 12406 10364 12434
rect 9680 12368 9732 12374
rect 9678 12336 9680 12345
rect 9732 12336 9734 12345
rect 9784 12306 9812 12406
rect 9678 12271 9734 12280
rect 9772 12300 9824 12306
rect 9692 11898 9720 12271
rect 9772 12242 9824 12248
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 9508 11342 9628 11370
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 8944 11076 8996 11082
rect 8944 11018 8996 11024
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 7944 4146 7972 8774
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 1216 3664 1268 3670
rect 1216 3606 1268 3612
rect 1228 400 1256 3606
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 3712 400 3740 4082
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 6196 400 6224 3674
rect 8404 3670 8432 7210
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 8588 2774 8616 8502
rect 8864 8430 8892 9590
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8956 6866 8984 11018
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9232 9042 9260 9318
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 9048 6730 9076 7278
rect 9324 6866 9352 11018
rect 9508 9654 9536 11342
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 10606 9628 11154
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9600 10198 9628 10542
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9692 9722 9720 10406
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 9864 10192 9916 10198
rect 9862 10160 9864 10169
rect 9916 10160 9918 10169
rect 9862 10095 9918 10104
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9496 9648 9548 9654
rect 9772 9648 9824 9654
rect 9548 9596 9720 9602
rect 9496 9590 9720 9596
rect 9824 9596 9996 9602
rect 9772 9590 9996 9596
rect 9508 9574 9720 9590
rect 9784 9586 9996 9590
rect 9784 9580 10008 9586
rect 9784 9574 9956 9580
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9110 9444 9454
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9692 8650 9720 9574
rect 9956 9522 10008 9528
rect 10060 9450 10088 9930
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 10152 9382 10180 9862
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9600 8622 9720 8650
rect 9600 8022 9628 8622
rect 9876 8498 9904 8842
rect 9864 8492 9916 8498
rect 9692 8452 9864 8480
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9600 6866 9628 7958
rect 9692 7410 9720 8452
rect 9864 8434 9916 8440
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10244 8090 10272 11018
rect 10336 9586 10364 12406
rect 10428 11286 10456 17070
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10704 16454 10732 17002
rect 11244 16720 11296 16726
rect 11244 16662 11296 16668
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10704 14958 10732 16390
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10692 14952 10744 14958
rect 10692 14894 10744 14900
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12986 10548 13330
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10704 12918 10732 13262
rect 10796 13258 10824 14350
rect 11072 13870 11100 15982
rect 11256 15586 11284 16662
rect 11348 16250 11376 17274
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 11336 16244 11388 16250
rect 11336 16186 11388 16192
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15706 11376 15982
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11704 15632 11756 15638
rect 11256 15558 11376 15586
rect 11704 15574 11756 15580
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 10968 13320 11020 13326
rect 11072 13308 11100 13806
rect 11020 13280 11100 13308
rect 10968 13262 11020 13268
rect 10784 13252 10836 13258
rect 10784 13194 10836 13200
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10612 10606 10640 11494
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 10169 10640 10542
rect 10598 10160 10654 10169
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10508 10124 10560 10130
rect 10598 10095 10654 10104
rect 10508 10066 10560 10072
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10336 9042 10364 9318
rect 10428 9178 10456 10066
rect 10520 9382 10548 10066
rect 10704 10062 10732 12854
rect 10782 11792 10838 11801
rect 10782 11727 10838 11736
rect 10796 11694 10824 11727
rect 10980 11694 11008 13262
rect 11164 13190 11192 14418
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 13870 11284 14214
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11348 13716 11376 15558
rect 11716 15434 11744 15574
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11716 14958 11744 15370
rect 11808 15162 11836 15506
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11992 15026 12020 15846
rect 12360 15502 12388 15846
rect 12452 15570 12480 16118
rect 12544 15570 12572 16186
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11440 14074 11468 14282
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11256 13688 11376 13716
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12782 11192 13126
rect 11152 12776 11204 12782
rect 11072 12736 11152 12764
rect 11072 12306 11100 12736
rect 11152 12718 11204 12724
rect 11256 12434 11284 13688
rect 11532 13274 11560 14826
rect 12636 14550 12664 18566
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15706 12848 15846
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12912 14890 12940 15914
rect 13096 15502 13124 16050
rect 13084 15496 13136 15502
rect 13082 15464 13084 15473
rect 13136 15464 13138 15473
rect 13082 15399 13138 15408
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 13096 15026 13124 15302
rect 13188 15162 13216 16186
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13280 15502 13308 15982
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15638 13400 15846
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13464 15502 13492 15914
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 12992 14952 13044 14958
rect 13280 14906 13308 15438
rect 13452 15360 13504 15366
rect 13556 15348 13584 15846
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 15570 13676 15642
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13504 15320 13584 15348
rect 13636 15360 13688 15366
rect 13452 15302 13504 15308
rect 13636 15302 13688 15308
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13044 14900 13308 14906
rect 12992 14894 13308 14900
rect 12900 14884 12952 14890
rect 13004 14878 13308 14894
rect 12900 14826 12952 14832
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 13464 14482 13492 15030
rect 13648 14958 13676 15302
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14482 13584 14758
rect 13924 14618 13952 15506
rect 14108 14958 14136 15846
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11624 13394 11652 14214
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11532 13246 11652 13274
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11164 12406 11284 12434
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 10198 10824 10542
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10980 10130 11008 10678
rect 11164 10266 11192 12406
rect 11244 12368 11296 12374
rect 11244 12310 11296 12316
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10784 9920 10836 9926
rect 10784 9862 10836 9868
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 8022 10364 8978
rect 10612 8090 10640 9386
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 9416 6458 9444 6802
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 5778 9536 6598
rect 9692 5846 9720 7346
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 9956 6928 10008 6934
rect 9956 6870 10008 6876
rect 9968 6254 9996 6870
rect 10152 6322 10180 6938
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8680 3738 8708 5510
rect 9692 5370 9720 5782
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 10244 5166 10272 7686
rect 10612 7410 10640 8026
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10520 6866 10548 7142
rect 10612 7002 10640 7346
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10704 6866 10732 9658
rect 10796 9518 10824 9862
rect 10888 9518 10916 10066
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8362 10824 9318
rect 11256 9110 11284 12310
rect 11348 9994 11376 12786
rect 11624 12782 11652 13246
rect 12084 13190 12112 14350
rect 13464 14278 13492 14418
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 13464 13802 13492 14214
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13452 13796 13504 13802
rect 13452 13738 13504 13744
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 13728 13728 13780 13734
rect 13728 13670 13780 13676
rect 12636 13462 12664 13670
rect 12728 13462 12756 13670
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12084 12918 12112 13126
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11612 12776 11664 12782
rect 12164 12776 12216 12782
rect 11612 12718 11664 12724
rect 12084 12736 12164 12764
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 11440 12306 11468 12582
rect 11532 12306 11560 12718
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 12084 12238 12112 12736
rect 12544 12730 12572 13126
rect 12636 12782 12664 13398
rect 12728 12782 12756 13398
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12164 12718 12216 12724
rect 12452 12702 12572 12730
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12452 12646 12480 12702
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11440 11694 11468 12038
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 12084 11558 12112 12174
rect 12544 12170 12572 12582
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 12544 11898 12572 12106
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12636 11218 12664 12718
rect 12912 12434 12940 12786
rect 12820 12406 12940 12434
rect 13096 12434 13124 12922
rect 13556 12782 13584 13262
rect 13740 13190 13768 13670
rect 13924 13394 13952 13874
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13556 12434 13584 12718
rect 13096 12406 13308 12434
rect 13556 12406 13676 12434
rect 12820 11762 12848 12406
rect 13280 11830 13308 12406
rect 13648 12306 13676 12406
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12636 10674 12664 11154
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12728 10606 12756 11630
rect 12820 11540 12848 11698
rect 12992 11552 13044 11558
rect 12820 11512 12992 11540
rect 12992 11494 13044 11500
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 13096 10810 13124 11222
rect 13280 11218 13308 11766
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 11348 9178 11376 9930
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11244 9104 11296 9110
rect 11244 9046 11296 9052
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 10980 7342 11008 7958
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10980 6934 11008 7278
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10692 6724 10744 6730
rect 10796 6712 10824 6802
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10744 6684 10824 6712
rect 10692 6666 10744 6672
rect 10704 6322 10732 6666
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10980 6254 11008 6598
rect 11164 6390 11192 6734
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 10968 6248 11020 6254
rect 10874 6216 10930 6225
rect 10968 6190 11020 6196
rect 10874 6151 10876 6160
rect 10928 6151 10930 6160
rect 10876 6122 10928 6128
rect 11072 5846 11100 6326
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10980 5234 11008 5714
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 11256 5098 11284 6666
rect 11624 5098 11652 9862
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 13004 9586 13032 9930
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12992 9580 13044 9586
rect 12992 9522 13044 9528
rect 12256 9512 12308 9518
rect 12308 9460 12480 9466
rect 12256 9454 12480 9460
rect 12268 9438 12480 9454
rect 12452 8906 12480 9438
rect 12440 8900 12492 8906
rect 12440 8842 12492 8848
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11808 8634 11836 8774
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 12544 8498 12572 9522
rect 12900 9512 12952 9518
rect 13096 9466 13124 10746
rect 13280 10606 13308 11154
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13188 9518 13216 9658
rect 13280 9586 13308 10406
rect 13372 10198 13400 10406
rect 13464 10266 13492 11698
rect 13648 11694 13676 12242
rect 13832 11898 13860 12718
rect 13924 12374 13952 13330
rect 14016 12986 14044 13330
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14200 12850 14228 18566
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14384 14890 14412 15982
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 14462 15464 14518 15473
rect 14462 15399 14518 15408
rect 14476 15094 14504 15399
rect 14936 15162 14964 15982
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15120 15162 15148 15302
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14414 14412 14826
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14384 12782 14412 13670
rect 14476 12850 14504 15030
rect 14936 14822 14964 15098
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14752 13802 14780 14282
rect 14936 13870 14964 14418
rect 15120 14074 15148 14418
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14740 13796 14792 13802
rect 14740 13738 14792 13744
rect 14936 13734 14964 13806
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 15120 13530 15148 13738
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14936 11694 14964 12786
rect 15120 12714 15148 13466
rect 15212 13462 15240 18566
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 17512 18222 17540 18566
rect 17500 18216 17552 18222
rect 17500 18158 17552 18164
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 15856 17814 15884 18022
rect 16960 17814 16988 18022
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 16948 17808 17000 17814
rect 16948 17750 17000 17756
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 15706 15332 17614
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 17880 17066 17908 17478
rect 16764 17060 16816 17066
rect 16764 17002 16816 17008
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15304 15026 15332 15642
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15396 15026 15424 15302
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15304 13870 15332 14962
rect 16776 14958 16804 17002
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 19076 16017 19104 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 19062 16008 19118 16017
rect 19062 15943 19118 15952
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 16868 14600 16896 15098
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 14618 16988 14894
rect 17408 14884 17460 14890
rect 17408 14826 17460 14832
rect 17132 14816 17184 14822
rect 17132 14758 17184 14764
rect 16776 14572 16896 14600
rect 16948 14612 17000 14618
rect 16580 14476 16632 14482
rect 16580 14418 16632 14424
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16488 14340 16540 14346
rect 16488 14282 16540 14288
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13870 15516 14214
rect 16500 13954 16528 14282
rect 16592 14074 16620 14418
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16500 13926 16620 13954
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15304 12850 15332 13806
rect 16120 13184 16172 13190
rect 16120 13126 16172 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 14924 11688 14976 11694
rect 14924 11630 14976 11636
rect 15028 11558 15056 12038
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15200 11688 15252 11694
rect 15120 11636 15200 11642
rect 15120 11630 15252 11636
rect 15120 11614 15240 11630
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14200 11234 14228 11494
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 14200 11206 14320 11234
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13360 10192 13412 10198
rect 13360 10134 13412 10140
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12900 9454 12952 9460
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 8498 12664 9318
rect 12912 9178 12940 9454
rect 13004 9438 13124 9466
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 8922 13032 9438
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9042 13124 9318
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13004 8906 13124 8922
rect 13004 8900 13136 8906
rect 13004 8894 13084 8900
rect 13084 8842 13136 8848
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 11716 7342 11744 8434
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7886 12020 8230
rect 12176 8090 12204 8366
rect 12452 8090 12480 8366
rect 13096 8362 13124 8842
rect 13188 8634 13216 8978
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12544 7954 12572 8191
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 12820 7546 12848 7890
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12162 6896 12218 6905
rect 12728 6866 12756 7278
rect 13096 7274 13124 8298
rect 13280 8294 13308 8910
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13280 7750 13308 8230
rect 13372 8090 13400 10134
rect 13464 9674 13492 10202
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9926 13952 9998
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13464 9646 13584 9674
rect 13556 8974 13584 9646
rect 13820 9648 13872 9654
rect 13634 9616 13690 9625
rect 13820 9590 13872 9596
rect 13634 9551 13690 9560
rect 13648 9518 13676 9551
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 9178 13676 9318
rect 13740 9178 13768 9386
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13450 8800 13506 8809
rect 13450 8735 13506 8744
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13464 7954 13492 8735
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 7002 13216 7142
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12162 6831 12164 6840
rect 12216 6831 12218 6840
rect 12624 6860 12676 6866
rect 12164 6802 12216 6808
rect 12624 6802 12676 6808
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12636 6746 12664 6802
rect 13188 6798 13216 6938
rect 13464 6934 13492 7890
rect 13556 7002 13584 8910
rect 13740 8809 13768 8910
rect 13726 8800 13782 8809
rect 13726 8735 13782 8744
rect 13832 8634 13860 9590
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13648 7886 13676 8366
rect 13924 8362 13952 9862
rect 14016 8974 14044 10474
rect 14108 10130 14136 10542
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9586 14136 9862
rect 14200 9625 14228 11086
rect 14292 9654 14320 11206
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14280 9648 14332 9654
rect 14186 9616 14242 9625
rect 14096 9580 14148 9586
rect 14280 9590 14332 9596
rect 14186 9551 14188 9560
rect 14096 9522 14148 9528
rect 14240 9551 14242 9560
rect 14188 9522 14240 9528
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 9042 14228 9318
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13740 8265 13768 8298
rect 13726 8256 13782 8265
rect 13782 8214 13860 8242
rect 13726 8191 13782 8200
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13740 6866 13768 7686
rect 13832 7410 13860 8214
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13924 6905 13952 8298
rect 14016 7342 14044 8910
rect 14292 8650 14320 9590
rect 14384 9081 14412 10610
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14542 10299 14850 10308
rect 14936 10130 14964 10746
rect 15028 10674 15056 11494
rect 15120 11218 15148 11614
rect 15948 11558 15976 11834
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 15120 10010 15148 10474
rect 15212 10198 15240 10542
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15304 10130 15332 11494
rect 16132 10130 16160 13126
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16500 12434 16528 12650
rect 16408 12406 16528 12434
rect 16592 12434 16620 13926
rect 16684 12918 16712 14418
rect 16776 13852 16804 14572
rect 16948 14554 17000 14560
rect 17144 14482 17172 14758
rect 17420 14482 17448 14826
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 16948 13864 17000 13870
rect 16776 13824 16948 13852
rect 16948 13806 17000 13812
rect 16960 13394 16988 13806
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12434 16896 12582
rect 16592 12406 16712 12434
rect 16408 11762 16436 12406
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16408 11218 16436 11698
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16408 10606 16436 11154
rect 16500 10742 16528 11494
rect 16684 11150 16712 12406
rect 16776 12406 16896 12434
rect 16776 11694 16804 12406
rect 17328 12306 17356 14214
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 16764 11688 16816 11694
rect 17328 11642 17356 12242
rect 16764 11630 16816 11636
rect 17236 11614 17356 11642
rect 16672 11144 16724 11150
rect 16592 11092 16672 11098
rect 16592 11086 16724 11092
rect 16592 11070 16712 11086
rect 17236 11082 17264 11614
rect 17420 11286 17448 14418
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17512 13394 17540 13874
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 12646 17540 13330
rect 17500 12640 17552 12646
rect 17500 12582 17552 12588
rect 17512 12306 17540 12582
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17408 11280 17460 11286
rect 17408 11222 17460 11228
rect 17224 11076 17276 11082
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15120 9982 15240 10010
rect 15212 9654 15240 9982
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9722 15332 9930
rect 16132 9926 16160 10066
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 9110 14504 9386
rect 15028 9382 15056 9454
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14464 9104 14516 9110
rect 14370 9072 14426 9081
rect 14464 9046 14516 9052
rect 14370 9007 14372 9016
rect 14424 9007 14426 9016
rect 14740 9036 14792 9042
rect 14372 8978 14424 8984
rect 14740 8978 14792 8984
rect 14464 8968 14516 8974
rect 14752 8945 14780 8978
rect 14464 8910 14516 8916
rect 14738 8936 14794 8945
rect 14108 8622 14320 8650
rect 14108 8430 14136 8622
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13910 6896 13966 6905
rect 13728 6860 13780 6866
rect 13910 6831 13966 6840
rect 13728 6802 13780 6808
rect 13176 6792 13228 6798
rect 12636 6730 12756 6746
rect 13176 6734 13228 6740
rect 12532 6724 12584 6730
rect 12636 6724 12768 6730
rect 12636 6718 12716 6724
rect 12532 6666 12584 6672
rect 12716 6666 12768 6672
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 12544 6322 12572 6666
rect 13740 6662 13768 6802
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 13556 6254 13584 6598
rect 14016 6254 14044 7142
rect 14200 6254 14228 8502
rect 14476 8430 14504 8910
rect 14738 8871 14794 8880
rect 14752 8498 14780 8871
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 14936 8090 14964 8366
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14292 7206 14320 7482
rect 14476 7342 14504 7890
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14370 6896 14426 6905
rect 14370 6831 14372 6840
rect 14424 6831 14426 6840
rect 14372 6802 14424 6808
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6390 14504 6598
rect 14660 6458 14688 6938
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14464 6384 14516 6390
rect 14464 6326 14516 6332
rect 14936 6254 14964 7890
rect 15028 7886 15056 9318
rect 15106 9072 15162 9081
rect 15106 9007 15162 9016
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15028 6798 15056 7278
rect 15120 7274 15148 9007
rect 15304 8974 15332 9658
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15304 8838 15332 8910
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8430 15332 8774
rect 15396 8430 15424 8978
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15292 8424 15344 8430
rect 15292 8366 15344 8372
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15212 8022 15240 8366
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15304 7886 15332 8366
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15108 7268 15160 7274
rect 15108 7210 15160 7216
rect 15292 7268 15344 7274
rect 15292 7210 15344 7216
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 15120 6254 15148 7210
rect 15304 6866 15332 7210
rect 15396 6934 15424 8366
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15488 7750 15516 8298
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15580 7206 15608 8366
rect 15672 8090 15700 8366
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15488 6866 15516 7142
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15212 6390 15240 6734
rect 15488 6390 15516 6802
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15672 6322 15700 7686
rect 15764 7410 15792 9522
rect 15856 9518 15884 9590
rect 15844 9512 15896 9518
rect 15896 9472 15976 9500
rect 15844 9454 15896 9460
rect 15948 8634 15976 9472
rect 16040 9178 16068 9590
rect 16132 9382 16160 9862
rect 16500 9382 16528 10678
rect 16592 10606 16620 11070
rect 17224 11018 17276 11024
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 17236 10606 17264 11018
rect 17408 11008 17460 11014
rect 17408 10950 17460 10956
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17420 10130 17448 10950
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9518 16620 9998
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 16948 9648 17000 9654
rect 16948 9590 17000 9596
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16120 9376 16172 9382
rect 16488 9376 16540 9382
rect 16172 9336 16252 9364
rect 16120 9318 16172 9324
rect 16224 9178 16252 9336
rect 16488 9318 16540 9324
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16500 9042 16528 9318
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16028 9036 16080 9042
rect 16028 8978 16080 8984
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16040 8838 16068 8978
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16132 8838 16160 8910
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16120 8832 16172 8838
rect 16224 8809 16252 8842
rect 16304 8832 16356 8838
rect 16120 8774 16172 8780
rect 16210 8800 16266 8809
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15764 6322 15792 7346
rect 15856 7342 15884 8434
rect 15948 7886 15976 8570
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 15948 7478 15976 7822
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6458 15884 7142
rect 16040 7002 16068 8774
rect 16132 8430 16160 8774
rect 16304 8774 16356 8780
rect 16210 8735 16266 8744
rect 16316 8634 16344 8774
rect 16500 8634 16528 8978
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16592 8430 16620 9114
rect 16670 9072 16726 9081
rect 16960 9042 16988 9590
rect 17420 9042 17448 10066
rect 17696 9586 17724 13942
rect 18156 13530 18184 14214
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18616 12986 18644 13262
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18420 12980 18472 12986
rect 18420 12922 18472 12928
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17880 10062 17908 11222
rect 18052 10532 18104 10538
rect 18052 10474 18104 10480
rect 18064 10266 18092 10474
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 9178 17724 9522
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 16670 9007 16726 9016
rect 16948 9036 17000 9042
rect 16684 8974 16712 9007
rect 16948 8978 17000 8984
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16592 7342 16620 8366
rect 16684 7993 16712 8910
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16670 7984 16726 7993
rect 17052 7954 17080 8502
rect 17420 8430 17448 8978
rect 17512 8945 17540 9114
rect 17696 9042 17724 9114
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17880 9024 17908 9998
rect 18064 9110 18092 10202
rect 18432 9897 18460 12922
rect 18800 12782 18828 13126
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 18418 9888 18474 9897
rect 18418 9823 18474 9832
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18052 9104 18104 9110
rect 18052 9046 18104 9052
rect 18248 9042 18276 9114
rect 17960 9036 18012 9042
rect 17880 8996 17960 9024
rect 17498 8936 17554 8945
rect 17498 8871 17554 8880
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17328 7954 17356 8298
rect 17512 8294 17540 8502
rect 17788 8498 17816 8978
rect 17880 8566 17908 8996
rect 17960 8978 18012 8984
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17500 8288 17552 8294
rect 17420 8248 17500 8276
rect 16670 7919 16726 7928
rect 17040 7948 17092 7954
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15844 6452 15896 6458
rect 15844 6394 15896 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 16592 6254 16620 7278
rect 16684 6934 16712 7919
rect 17040 7890 17092 7896
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17236 7342 17264 7482
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16868 6662 16896 7142
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 17236 6254 17264 7278
rect 17420 7206 17448 8248
rect 17500 8230 17552 8236
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17498 7984 17554 7993
rect 17604 7954 17632 8230
rect 17972 7954 18000 8842
rect 18248 8294 18276 8978
rect 18432 8430 18460 8978
rect 18420 8424 18472 8430
rect 18420 8366 18472 8372
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 17498 7919 17500 7928
rect 17552 7919 17554 7928
rect 17592 7948 17644 7954
rect 17500 7890 17552 7896
rect 17592 7890 17644 7896
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17512 7410 17540 7686
rect 18064 7546 18092 7686
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 7200 17460 7206
rect 17408 7142 17460 7148
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 6458 17356 6598
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17328 6254 17356 6394
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 16580 6248 16632 6254
rect 16948 6248 17000 6254
rect 16580 6190 16632 6196
rect 16776 6196 16948 6202
rect 16776 6190 17000 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 16776 6186 16988 6190
rect 16764 6180 16988 6186
rect 16816 6174 16988 6180
rect 16764 6122 16816 6128
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11060 5024 11112 5030
rect 11060 4966 11112 4972
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8588 2746 8708 2774
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 8680 400 8708 2746
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 11072 2530 11100 4966
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 11072 2502 11192 2530
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 11164 400 11192 2502
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 13648 400 13676 5510
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 16132 400 16160 4966
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 18616 400 18644 4966
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
rect 11150 0 11206 400
rect 13634 0 13690 400
rect 16118 0 16174 400
rect 18602 0 18658 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 7102 12552 7158 12608
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 10322 16632 10378 16688
rect 9678 12316 9680 12336
rect 9680 12316 9732 12336
rect 9732 12316 9734 12336
rect 9678 12280 9734 12316
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 9862 10140 9864 10160
rect 9864 10140 9916 10160
rect 9916 10140 9918 10160
rect 9862 10104 9918 10140
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 10598 10104 10654 10160
rect 10782 11736 10838 11792
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 13082 15444 13084 15464
rect 13084 15444 13136 15464
rect 13136 15444 13138 15464
rect 13082 15408 13138 15444
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 10874 6180 10930 6216
rect 10874 6160 10876 6180
rect 10876 6160 10928 6180
rect 10928 6160 10930 6180
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 14462 15408 14518 15464
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 19062 15952 19118 16008
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 12530 8200 12586 8256
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 12162 6860 12218 6896
rect 13634 9560 13690 9616
rect 13450 8744 13506 8800
rect 12162 6840 12164 6860
rect 12164 6840 12216 6860
rect 12216 6840 12218 6860
rect 13726 8744 13782 8800
rect 14186 9580 14242 9616
rect 14186 9560 14188 9580
rect 14188 9560 14240 9580
rect 14240 9560 14242 9580
rect 13726 8200 13782 8256
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 14370 9036 14426 9072
rect 14370 9016 14372 9036
rect 14372 9016 14424 9036
rect 14424 9016 14426 9036
rect 13910 6840 13966 6896
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 14738 8880 14794 8936
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 14370 6860 14426 6896
rect 14370 6840 14372 6860
rect 14372 6840 14424 6860
rect 14424 6840 14426 6860
rect 15106 9016 15162 9072
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 16210 8744 16266 8800
rect 16670 9016 16726 9072
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 16670 7928 16726 7984
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 18418 9832 18474 9888
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 17498 8880 17554 8936
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17498 7948 17554 7984
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 17498 7928 17500 7948
rect 17500 7928 17552 7948
rect 17552 7928 17554 7948
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 10317 16690 10383 16693
rect 10910 16690 10916 16692
rect 10317 16688 10916 16690
rect 10317 16632 10322 16688
rect 10378 16632 10916 16688
rect 10317 16630 10916 16632
rect 10317 16627 10383 16630
rect 10910 16628 10916 16630
rect 10980 16628 10986 16692
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 19057 16010 19123 16013
rect 17972 16008 19123 16010
rect 17972 15952 19062 16008
rect 19118 15952 19123 16008
rect 17972 15950 19123 15952
rect 17972 15948 17978 15950
rect 19057 15947 19123 15950
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 13077 15466 13143 15469
rect 14457 15466 14523 15469
rect 13077 15464 14523 15466
rect 13077 15408 13082 15464
rect 13138 15408 14462 15464
rect 14518 15408 14523 15464
rect 13077 15406 14523 15408
rect 13077 15403 13143 15406
rect 14457 15403 14523 15406
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 7097 12610 7163 12613
rect 7097 12608 7298 12610
rect 7097 12552 7102 12608
rect 7158 12552 7298 12608
rect 7097 12550 7298 12552
rect 7097 12547 7163 12550
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 7238 12338 7298 12550
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 9673 12338 9739 12341
rect 7238 12336 9739 12338
rect 7238 12280 9678 12336
rect 9734 12280 9739 12336
rect 7238 12278 9739 12280
rect 9673 12275 9739 12278
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 10777 11794 10843 11797
rect 17902 11794 17908 11796
rect 10777 11792 17908 11794
rect 10777 11736 10782 11792
rect 10838 11736 17908 11792
rect 10777 11734 17908 11736
rect 10777 11731 10843 11734
rect 17902 11732 17908 11734
rect 17972 11732 17978 11796
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 9857 10162 9923 10165
rect 10593 10162 10659 10165
rect 9857 10160 10659 10162
rect 9857 10104 9862 10160
rect 9918 10104 10598 10160
rect 10654 10104 10659 10160
rect 9857 10102 10659 10104
rect 9857 10099 9923 10102
rect 10593 10099 10659 10102
rect 18413 9890 18479 9893
rect 19600 9890 20000 9920
rect 18413 9888 20000 9890
rect 18413 9832 18418 9888
rect 18474 9832 20000 9888
rect 18413 9830 20000 9832
rect 18413 9827 18479 9830
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 19600 9800 20000 9830
rect 16896 9759 17212 9760
rect 13629 9618 13695 9621
rect 14181 9618 14247 9621
rect 13629 9616 14247 9618
rect 13629 9560 13634 9616
rect 13690 9560 14186 9616
rect 14242 9560 14247 9616
rect 13629 9558 14247 9560
rect 13629 9555 13695 9558
rect 14181 9555 14247 9558
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 14365 9074 14431 9077
rect 15101 9074 15167 9077
rect 16665 9074 16731 9077
rect 14365 9072 16731 9074
rect 14365 9016 14370 9072
rect 14426 9016 15106 9072
rect 15162 9016 16670 9072
rect 16726 9016 16731 9072
rect 14365 9014 16731 9016
rect 14365 9011 14431 9014
rect 15101 9011 15167 9014
rect 16665 9011 16731 9014
rect 14733 8938 14799 8941
rect 17493 8938 17559 8941
rect 14733 8936 17559 8938
rect 14733 8880 14738 8936
rect 14794 8880 17498 8936
rect 17554 8880 17559 8936
rect 14733 8878 17559 8880
rect 14733 8875 14799 8878
rect 17493 8875 17559 8878
rect 13445 8802 13511 8805
rect 13721 8802 13787 8805
rect 16205 8802 16271 8805
rect 13445 8800 16271 8802
rect 13445 8744 13450 8800
rect 13506 8744 13726 8800
rect 13782 8744 16210 8800
rect 16266 8744 16271 8800
rect 13445 8742 16271 8744
rect 13445 8739 13511 8742
rect 13721 8739 13787 8742
rect 16205 8739 16271 8742
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 12525 8258 12591 8261
rect 13721 8258 13787 8261
rect 12525 8256 13787 8258
rect 12525 8200 12530 8256
rect 12586 8200 13726 8256
rect 13782 8200 13787 8256
rect 12525 8198 13787 8200
rect 12525 8195 12591 8198
rect 13721 8195 13787 8198
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19253 8127 19569 8128
rect 16665 7986 16731 7989
rect 17493 7986 17559 7989
rect 16665 7984 17559 7986
rect 16665 7928 16670 7984
rect 16726 7928 17498 7984
rect 17554 7928 17559 7984
rect 16665 7926 17559 7928
rect 16665 7923 16731 7926
rect 17493 7923 17559 7926
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 12157 6898 12223 6901
rect 13905 6898 13971 6901
rect 14365 6898 14431 6901
rect 12157 6896 14431 6898
rect 12157 6840 12162 6896
rect 12218 6840 13910 6896
rect 13966 6840 14370 6896
rect 14426 6840 14431 6896
rect 12157 6838 14431 6840
rect 12157 6835 12223 6838
rect 13905 6835 13971 6838
rect 14365 6835 14431 6838
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 10869 6220 10935 6221
rect 10869 6218 10916 6220
rect 10824 6216 10916 6218
rect 10824 6160 10874 6216
rect 10824 6158 10916 6160
rect 10869 6156 10916 6158
rect 10980 6156 10986 6220
rect 10869 6155 10935 6156
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 10916 16628 10980 16692
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 17908 15948 17972 16012
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 17908 11732 17972 11796
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 10916 6216 10980 6220
rect 10916 6160 10930 6216
rect 10930 6160 10980 6216
rect 10916 6156 10980 6160
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 10918 6221 10978 16627
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 10915 6220 10981 6221
rect 10915 6156 10916 6220
rect 10980 6156 10981 6220
rect 10915 6155 10981 6156
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 17907 16012 17973 16013
rect 17907 15948 17908 16012
rect 17972 15948 17973 16012
rect 17907 15947 17973 15948
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 17910 11797 17970 15947
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 17907 11796 17973 11797
rect 17907 11732 17908 11796
rect 17972 11732 17973 11796
rect 17907 11731 17973 11732
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__inv_2  _214_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 1704896540
transform -1 0 8924 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 1704896540
transform -1 0 8188 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1704896540
transform 1 0 5980 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _218_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7268 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1704896540
transform 1 0 6716 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 1704896540
transform 1 0 6256 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6256 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _224_
timestamp 1704896540
transform 1 0 6992 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _225_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6992 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _228_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6808 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _232_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11960 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11224 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4508 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _237_
timestamp 1704896540
transform -1 0 5612 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp 1704896540
transform -1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4692 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp 1704896540
transform -1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _241_
timestamp 1704896540
transform -1 0 4508 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1704896540
transform 1 0 3956 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5152 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp 1704896540
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _245_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6072 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _246_
timestamp 1704896540
transform 1 0 5152 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _247_
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1704896540
transform -1 0 6716 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _249_
timestamp 1704896540
transform -1 0 5428 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4508 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _251_
timestamp 1704896540
transform 1 0 4508 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _252_
timestamp 1704896540
transform -1 0 4968 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _253_
timestamp 1704896540
transform -1 0 4784 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _254_
timestamp 1704896540
transform -1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _255_
timestamp 1704896540
transform -1 0 3680 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _256_
timestamp 1704896540
transform -1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _257_
timestamp 1704896540
transform -1 0 2576 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _259_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3772 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _260_
timestamp 1704896540
transform -1 0 3128 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2576 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _262_
timestamp 1704896540
transform 1 0 2024 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _263_
timestamp 1704896540
transform 1 0 2024 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _264_
timestamp 1704896540
transform -1 0 1932 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _265_
timestamp 1704896540
transform -1 0 1472 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _266_
timestamp 1704896540
transform -1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp 1704896540
transform 1 0 2392 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _268_
timestamp 1704896540
transform -1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _269_
timestamp 1704896540
transform 1 0 2668 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp 1704896540
transform -1 0 3036 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _271_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3956 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _272_
timestamp 1704896540
transform 1 0 8740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1704896540
transform 1 0 10028 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10948 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15456 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15916 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _278_
timestamp 1704896540
transform -1 0 12788 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _279_
timestamp 1704896540
transform 1 0 14352 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _280_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12788 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _281_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11868 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 18492 0 -1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _283_
timestamp 1704896540
transform 1 0 17020 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_2  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17848 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _285_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16376 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _286_
timestamp 1704896540
transform 1 0 16376 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _287_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 17020 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _288_
timestamp 1704896540
transform 1 0 14996 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _289_
timestamp 1704896540
transform -1 0 18124 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _290_
timestamp 1704896540
transform -1 0 16928 0 1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _291_
timestamp 1704896540
transform 1 0 15824 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _292_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12236 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _293_
timestamp 1704896540
transform -1 0 17112 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _294_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _295_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17480 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _296_
timestamp 1704896540
transform 1 0 15272 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _297_
timestamp 1704896540
transform 1 0 15088 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _298_
timestamp 1704896540
transform 1 0 16928 0 1 10336
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _299_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16560 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _300_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _301_
timestamp 1704896540
transform 1 0 17572 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _302_
timestamp 1704896540
transform 1 0 18032 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _303_
timestamp 1704896540
transform 1 0 17020 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _304_
timestamp 1704896540
transform -1 0 13800 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _305_
timestamp 1704896540
transform 1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _306_
timestamp 1704896540
transform 1 0 15180 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _307_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14444 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1704896540
transform 1 0 9568 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _309_
timestamp 1704896540
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _310_
timestamp 1704896540
transform 1 0 9752 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _311_
timestamp 1704896540
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _312_
timestamp 1704896540
transform 1 0 15824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _313_
timestamp 1704896540
transform 1 0 13800 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _314_
timestamp 1704896540
transform -1 0 13984 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _315_
timestamp 1704896540
transform -1 0 13156 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _316_
timestamp 1704896540
transform 1 0 18216 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _317_
timestamp 1704896540
transform -1 0 15180 0 -1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _318_
timestamp 1704896540
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _319_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16928 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _320_
timestamp 1704896540
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _321_
timestamp 1704896540
transform -1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _322_
timestamp 1704896540
transform 1 0 15456 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _323_
timestamp 1704896540
transform -1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _324_
timestamp 1704896540
transform 1 0 12880 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _325_
timestamp 1704896540
transform 1 0 11868 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp 1704896540
transform 1 0 10580 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _327_
timestamp 1704896540
transform 1 0 10028 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _328_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _329_
timestamp 1704896540
transform 1 0 10672 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _330_
timestamp 1704896540
transform 1 0 9200 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _331_
timestamp 1704896540
transform 1 0 9108 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _332_
timestamp 1704896540
transform 1 0 16192 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _333_
timestamp 1704896540
transform 1 0 16652 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _334_
timestamp 1704896540
transform 1 0 17204 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _335_
timestamp 1704896540
transform 1 0 16836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _336_
timestamp 1704896540
transform 1 0 14444 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _337_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14720 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _338_
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _339_
timestamp 1704896540
transform -1 0 14720 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _340_
timestamp 1704896540
transform 1 0 14076 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _341_
timestamp 1704896540
transform 1 0 16284 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _342_
timestamp 1704896540
transform 1 0 14352 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _343_
timestamp 1704896540
transform -1 0 14536 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _344_
timestamp 1704896540
transform 1 0 13708 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp 1704896540
transform -1 0 14444 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _346_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13524 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _347_
timestamp 1704896540
transform 1 0 13800 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _348_
timestamp 1704896540
transform 1 0 9660 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _349_
timestamp 1704896540
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _350_
timestamp 1704896540
transform -1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _351_
timestamp 1704896540
transform -1 0 18216 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _352_
timestamp 1704896540
transform -1 0 14628 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _353_
timestamp 1704896540
transform 1 0 13616 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _354_
timestamp 1704896540
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_1  _355_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15364 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _356_
timestamp 1704896540
transform 1 0 14168 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _357_
timestamp 1704896540
transform 1 0 14996 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _358_
timestamp 1704896540
transform 1 0 14812 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _359_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14076 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _360_
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1704896540
transform 1 0 9752 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _362_
timestamp 1704896540
transform 1 0 8832 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp 1704896540
transform -1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _364_
timestamp 1704896540
transform -1 0 13156 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _365_
timestamp 1704896540
transform 1 0 12880 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _366_
timestamp 1704896540
transform 1 0 12236 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _367_
timestamp 1704896540
transform 1 0 12144 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _368_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11960 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _370_
timestamp 1704896540
transform 1 0 9752 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _371_
timestamp 1704896540
transform -1 0 10488 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _373_
timestamp 1704896540
transform 1 0 11960 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _374_
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _375_
timestamp 1704896540
transform -1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _376_
timestamp 1704896540
transform -1 0 8648 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _377_
timestamp 1704896540
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _378_
timestamp 1704896540
transform -1 0 10856 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _379_
timestamp 1704896540
transform -1 0 11684 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _380_
timestamp 1704896540
transform -1 0 17112 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _381_
timestamp 1704896540
transform 1 0 12052 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11316 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _383_
timestamp 1704896540
transform 1 0 12788 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _384_
timestamp 1704896540
transform -1 0 14628 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _385_
timestamp 1704896540
transform -1 0 12972 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _386_
timestamp 1704896540
transform 1 0 12972 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1704896540
transform -1 0 15456 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _388_
timestamp 1704896540
transform 1 0 13524 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _389_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13892 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _390_
timestamp 1704896540
transform -1 0 13616 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _391_
timestamp 1704896540
transform -1 0 13800 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _392_
timestamp 1704896540
transform -1 0 13616 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _393_
timestamp 1704896540
transform -1 0 15180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _394_
timestamp 1704896540
transform -1 0 15548 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _395_
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _396_
timestamp 1704896540
transform 1 0 12512 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _397_
timestamp 1704896540
transform 1 0 12972 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _398_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11592 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _399_
timestamp 1704896540
transform 1 0 10948 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _400_
timestamp 1704896540
transform 1 0 10304 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _401_
timestamp 1704896540
transform -1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _402_
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _403_
timestamp 1704896540
transform 1 0 12052 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _404_
timestamp 1704896540
transform -1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _405_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11040 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _406_
timestamp 1704896540
transform 1 0 16836 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _407_
timestamp 1704896540
transform 1 0 12788 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _408_
timestamp 1704896540
transform 1 0 16928 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _409_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18124 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _410_
timestamp 1704896540
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _411_
timestamp 1704896540
transform 1 0 7636 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _412_
timestamp 1704896540
transform 1 0 8096 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _413_
timestamp 1704896540
transform 1 0 9016 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _414_
timestamp 1704896540
transform -1 0 9568 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _415_
timestamp 1704896540
transform 1 0 8648 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _416_
timestamp 1704896540
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _417_
timestamp 1704896540
transform 1 0 8924 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _418_
timestamp 1704896540
transform 1 0 9476 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _419_
timestamp 1704896540
transform -1 0 10120 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _420_
timestamp 1704896540
transform -1 0 9936 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _421_
timestamp 1704896540
transform 1 0 7728 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _422_
timestamp 1704896540
transform 1 0 8188 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _423_
timestamp 1704896540
transform 1 0 6532 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _424_
timestamp 1704896540
transform 1 0 6992 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _425_
timestamp 1704896540
transform -1 0 7728 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _426_
timestamp 1704896540
transform -1 0 7636 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _427_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp 1704896540
transform -1 0 6532 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp 1704896540
transform 1 0 3956 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp 1704896540
transform 1 0 6348 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp 1704896540
transform 1 0 4140 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _432_
timestamp 1704896540
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp 1704896540
transform 1 0 2024 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp 1704896540
transform -1 0 2300 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _435_
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _436_
timestamp 1704896540
transform -1 0 2300 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _437_
timestamp 1704896540
transform -1 0 3128 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _438_
timestamp 1704896540
transform 1 0 2024 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _439_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10120 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _440_
timestamp 1704896540
transform -1 0 9568 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _441_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10120 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _442_
timestamp 1704896540
transform -1 0 9936 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _443_
timestamp 1704896540
transform 1 0 9384 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _444_
timestamp 1704896540
transform 1 0 11316 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _445_
timestamp 1704896540
transform 1 0 10948 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _446_
timestamp 1704896540
transform 1 0 16652 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _447__12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15916 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _447_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 16100 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_4  _448_
timestamp 1704896540
transform 1 0 11040 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _449_
timestamp 1704896540
transform 1 0 15088 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _450_
timestamp 1704896540
transform 1 0 13616 0 -1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp 1704896540
transform 1 0 15180 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _452_
timestamp 1704896540
transform 1 0 11132 0 1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp 1704896540
transform 1 0 13892 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp 1704896540
transform 1 0 10856 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _456_
timestamp 1704896540
transform 1 0 17020 0 1 12512
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp 1704896540
transform -1 0 9016 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp 1704896540
transform 1 0 8464 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp 1704896540
transform -1 0 10028 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _460_
timestamp 1704896540
transform 1 0 9384 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _461_
timestamp 1704896540
transform 1 0 9108 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _462_
timestamp 1704896540
transform 1 0 8372 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _463_
timestamp 1704896540
transform -1 0 7268 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _464_
timestamp 1704896540
transform 1 0 4324 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10856 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 7176 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform -1 0 8280 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 11040 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 12328 0 -1 12512
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1704896540
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_201
timestamp 1704896540
transform 1 0 19044 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_193 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 18308 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp 1704896540
transform 1 0 19044 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1704896540
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1704896540
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 1704896540
transform 1 0 18676 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 1704896540
transform 1 0 19044 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_193
timestamp 1704896540
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 1704896540
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1704896540
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1704896540
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp 1704896540
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp 1704896540
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1704896540
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp 1704896540
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1704896540
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1704896540
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1704896540
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1704896540
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp 1704896540
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_201
timestamp 1704896540
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1704896540
transform 1 0 9108 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_130
timestamp 1704896540
transform 1 0 12512 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_165
timestamp 1704896540
transform 1 0 15732 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_173
timestamp 1704896540
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_192
timestamp 1704896540
transform 1 0 18216 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_197
timestamp 1704896540
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_201
timestamp 1704896540
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8004 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1704896540
transform 1 0 10120 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_134
timestamp 1704896540
transform 1 0 12880 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_146
timestamp 1704896540
transform 1 0 13984 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_158
timestamp 1704896540
transform 1 0 15088 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16100 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17204 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_193
timestamp 1704896540
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_201
timestamp 1704896540
transform 1 0 19044 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_97
timestamp 1704896540
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_108
timestamp 1704896540
transform 1 0 10488 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_115
timestamp 1704896540
transform 1 0 11132 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_127
timestamp 1704896540
transform 1 0 12236 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_151
timestamp 1704896540
transform 1 0 14444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_165
timestamp 1704896540
transform 1 0 15732 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_169
timestamp 1704896540
transform 1 0 16100 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_185
timestamp 1704896540
transform 1 0 17572 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1704896540
transform 1 0 18308 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1704896540
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1704896540
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8004 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_97
timestamp 1704896540
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_107
timestamp 1704896540
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_122
timestamp 1704896540
transform 1 0 11776 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_139
timestamp 1704896540
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1704896540
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16100 0 -1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_180
timestamp 1704896540
transform 1 0 17112 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_192
timestamp 1704896540
transform 1 0 18216 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_200
timestamp 1704896540
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_104
timestamp 1704896540
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_108
timestamp 1704896540
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_118
timestamp 1704896540
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_126
timestamp 1704896540
transform 1 0 12144 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_152
timestamp 1704896540
transform 1 0 14536 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_156
timestamp 1704896540
transform 1 0 14904 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_162
timestamp 1704896540
transform 1 0 15456 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_172
timestamp 1704896540
transform 1 0 16376 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_178
timestamp 1704896540
transform 1 0 16928 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_185
timestamp 1704896540
transform 1 0 17572 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1704896540
transform 1 0 18308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1704896540
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1704896540
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9108 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_99
timestamp 1704896540
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_104
timestamp 1704896540
transform 1 0 10120 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_122
timestamp 1704896540
transform 1 0 11776 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_144
timestamp 1704896540
transform 1 0 13800 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_150
timestamp 1704896540
transform 1 0 14352 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_154
timestamp 1704896540
transform 1 0 14720 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1704896540
transform 1 0 15732 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16100 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_177
timestamp 1704896540
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_193
timestamp 1704896540
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_201
timestamp 1704896540
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_102
timestamp 1704896540
transform 1 0 9936 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_114
timestamp 1704896540
transform 1 0 11040 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_137
timestamp 1704896540
transform 1 0 13156 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_168
timestamp 1704896540
transform 1 0 16008 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1704896540
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1704896540
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1704896540
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_77
timestamp 1704896540
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_98
timestamp 1704896540
transform 1 0 9568 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_102
timestamp 1704896540
transform 1 0 9936 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_106
timestamp 1704896540
transform 1 0 10304 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_141
timestamp 1704896540
transform 1 0 13524 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_157
timestamp 1704896540
transform 1 0 14996 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_161
timestamp 1704896540
transform 1 0 15364 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_195
timestamp 1704896540
transform 1 0 18492 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_201
timestamp 1704896540
transform 1 0 19044 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1704896540
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 1704896540
transform 1 0 8740 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_113
timestamp 1704896540
transform 1 0 10948 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_121
timestamp 1704896540
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1704896540
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_165
timestamp 1704896540
transform 1 0 15732 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_169
timestamp 1704896540
transform 1 0 16100 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_181
timestamp 1704896540
transform 1 0 17204 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1704896540
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 1704896540
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp 1704896540
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1704896540
transform 1 0 6900 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1704896540
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9108 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_121
timestamp 1704896540
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_133
timestamp 1704896540
transform 1 0 12788 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_141
timestamp 1704896540
transform 1 0 13524 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1704896540
transform 1 0 15364 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_177
timestamp 1704896540
transform 1 0 16836 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_184
timestamp 1704896540
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_196
timestamp 1704896540
transform 1 0 18584 0 -1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1704896540
transform 1 0 6532 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1704896540
transform 1 0 7636 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_88
timestamp 1704896540
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_100
timestamp 1704896540
transform 1 0 9752 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_106
timestamp 1704896540
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_113
timestamp 1704896540
transform 1 0 10948 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_125
timestamp 1704896540
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_191
timestamp 1704896540
transform 1 0 18124 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1704896540
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1704896540
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1704896540
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_32
timestamp 1704896540
transform 1 0 3496 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_60
timestamp 1704896540
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_72
timestamp 1704896540
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_84
timestamp 1704896540
transform 1 0 8280 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_88
timestamp 1704896540
transform 1 0 8648 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_92
timestamp 1704896540
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 1704896540
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1704896540
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 1704896540
transform 1 0 13892 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_159
timestamp 1704896540
transform 1 0 15180 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp 1704896540
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_65
timestamp 1704896540
transform 1 0 6532 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_71
timestamp 1704896540
transform 1 0 7084 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1704896540
transform 1 0 8924 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1704896540
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_153
timestamp 1704896540
transform 1 0 14628 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_162
timestamp 1704896540
transform 1 0 15456 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_166
timestamp 1704896540
transform 1 0 15824 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_180
timestamp 1704896540
transform 1 0 17112 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1704896540
transform 1 0 18216 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1704896540
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1704896540
transform 1 0 19044 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_19
timestamp 1704896540
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_25
timestamp 1704896540
transform 1 0 2852 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_43
timestamp 1704896540
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 5612 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1704896540
transform 1 0 6164 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_75
timestamp 1704896540
transform 1 0 7452 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_99
timestamp 1704896540
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_119
timestamp 1704896540
transform 1 0 11500 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_148
timestamp 1704896540
transform 1 0 14168 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_160
timestamp 1704896540
transform 1 0 15272 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_195
timestamp 1704896540
transform 1 0 18492 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp 1704896540
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_35
timestamp 1704896540
transform 1 0 3772 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_47
timestamp 1704896540
transform 1 0 4876 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_51
timestamp 1704896540
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_72
timestamp 1704896540
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_76
timestamp 1704896540
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_102
timestamp 1704896540
transform 1 0 9936 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_110
timestamp 1704896540
transform 1 0 10672 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_117
timestamp 1704896540
transform 1 0 11316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_123
timestamp 1704896540
transform 1 0 11868 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_147
timestamp 1704896540
transform 1 0 14076 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_155
timestamp 1704896540
transform 1 0 14812 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1704896540
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1704896540
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_23
timestamp 1704896540
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_33
timestamp 1704896540
transform 1 0 3588 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_41
timestamp 1704896540
transform 1 0 4324 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_45
timestamp 1704896540
transform 1 0 4692 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1704896540
transform 1 0 5428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_65
timestamp 1704896540
transform 1 0 6532 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_70
timestamp 1704896540
transform 1 0 6992 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_98
timestamp 1704896540
transform 1 0 9568 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_104
timestamp 1704896540
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1704896540
transform 1 0 12420 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_199
timestamp 1704896540
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1704896540
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_60
timestamp 1704896540
transform 1 0 6072 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1704896540
transform 1 0 7820 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8188 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1704896540
transform 1 0 9476 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_109
timestamp 1704896540
transform 1 0 10580 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_145
timestamp 1704896540
transform 1 0 13892 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_153
timestamp 1704896540
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_188
timestamp 1704896540
transform 1 0 17848 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp 1704896540
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_201
timestamp 1704896540
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_31
timestamp 1704896540
transform 1 0 3404 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 5612 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_79
timestamp 1704896540
transform 1 0 7820 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_83
timestamp 1704896540
transform 1 0 8188 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_89
timestamp 1704896540
transform 1 0 8740 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_98
timestamp 1704896540
transform 1 0 9568 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1704896540
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_113
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_128
timestamp 1704896540
transform 1 0 12328 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_136
timestamp 1704896540
transform 1 0 13064 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_142
timestamp 1704896540
transform 1 0 13616 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_154
timestamp 1704896540
transform 1 0 14720 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_163
timestamp 1704896540
transform 1 0 15548 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 15916 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16100 0 -1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_184
timestamp 1704896540
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_196
timestamp 1704896540
transform 1 0 18584 0 -1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_15
timestamp 1704896540
transform 1 0 1932 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4324 0 1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_51
timestamp 1704896540
transform 1 0 5244 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_63
timestamp 1704896540
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_103
timestamp 1704896540
transform 1 0 10028 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_109
timestamp 1704896540
transform 1 0 10580 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_116
timestamp 1704896540
transform 1 0 11224 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_124
timestamp 1704896540
transform 1 0 11960 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_132
timestamp 1704896540
transform 1 0 12696 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_144
timestamp 1704896540
transform 1 0 13800 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_155
timestamp 1704896540
transform 1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_182
timestamp 1704896540
transform 1 0 17296 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1704896540
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1704896540
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp 1704896540
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_19
timestamp 1704896540
transform 1 0 2300 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_35
timestamp 1704896540
transform 1 0 3772 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_46
timestamp 1704896540
transform 1 0 4784 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1704896540
transform 1 0 5520 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_57
timestamp 1704896540
transform 1 0 5796 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_65
timestamp 1704896540
transform 1 0 6532 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_93
timestamp 1704896540
transform 1 0 9108 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_102
timestamp 1704896540
transform 1 0 9936 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1704896540
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1704896540
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_162
timestamp 1704896540
transform 1 0 15456 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_193
timestamp 1704896540
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_201
timestamp 1704896540
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_3
timestamp 1704896540
transform 1 0 828 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 1704896540
transform 1 0 2668 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_42
timestamp 1704896540
transform 1 0 4416 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_53
timestamp 1704896540
transform 1 0 5428 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_61
timestamp 1704896540
transform 1 0 6164 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_67
timestamp 1704896540
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1704896540
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8372 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_109
timestamp 1704896540
transform 1 0 10580 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_113
timestamp 1704896540
transform 1 0 10948 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_133
timestamp 1704896540
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1704896540
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1704896540
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1704896540
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1704896540
transform 1 0 17940 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1704896540
transform 1 0 18492 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1704896540
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1704896540
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_15
timestamp 1704896540
transform 1 0 1932 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_32
timestamp 1704896540
transform 1 0 3496 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_38
timestamp 1704896540
transform 1 0 4048 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 5612 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_65
timestamp 1704896540
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_77
timestamp 1704896540
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_89
timestamp 1704896540
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_104
timestamp 1704896540
transform 1 0 10120 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1704896540
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1704896540
transform 1 0 12052 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1704896540
transform 1 0 13156 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1704896540
transform 1 0 14260 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1704896540
transform 1 0 15364 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 15916 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp 1704896540
transform 1 0 18308 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp 1704896540
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 828 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_15
timestamp 1704896540
transform 1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_22
timestamp 1704896540
transform 1 0 2576 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3220 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_35
timestamp 1704896540
transform 1 0 3772 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_39
timestamp 1704896540
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_46
timestamp 1704896540
transform 1 0 4784 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_58
timestamp 1704896540
transform 1 0 5888 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_65
timestamp 1704896540
transform 1 0 6532 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1704896540
transform 1 0 7636 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1704896540
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1704896540
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_91
timestamp 1704896540
transform 1 0 8924 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_108
timestamp 1704896540
transform 1 0 10488 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_114
timestamp 1704896540
transform 1 0 11040 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_119
timestamp 1704896540
transform 1 0 11500 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_131
timestamp 1704896540
transform 1 0 12604 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1704896540
transform 1 0 13340 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1704896540
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1704896540
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1704896540
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1704896540
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1704896540
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 1704896540
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp 1704896540
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1704896540
transform 1 0 828 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1704896540
transform 1 0 1932 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_27
timestamp 1704896540
transform 1 0 3036 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_35
timestamp 1704896540
transform 1 0 3772 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1704896540
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_116
timestamp 1704896540
transform 1 0 11224 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_128
timestamp 1704896540
transform 1 0 12328 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_140
timestamp 1704896540
transform 1 0 13432 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_152
timestamp 1704896540
transform 1 0 14536 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_164
timestamp 1704896540
transform 1 0 15640 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 1704896540
transform 1 0 18032 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1704896540
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1704896540
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1704896540
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1704896540
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_78
timestamp 1704896540
transform 1 0 7728 0 1 17952
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_108
timestamp 1704896540
transform 1 0 10488 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_120
timestamp 1704896540
transform 1 0 11592 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_132
timestamp 1704896540
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1704896540
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_153
timestamp 1704896540
transform 1 0 14628 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_161
timestamp 1704896540
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_167
timestamp 1704896540
transform 1 0 15916 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_175
timestamp 1704896540
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_180
timestamp 1704896540
transform 1 0 17112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1704896540
transform 1 0 18216 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1704896540
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp 1704896540
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1704896540
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_14
timestamp 1704896540
transform 1 0 1840 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp 1704896540
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_29
timestamp 1704896540
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_37
timestamp 1704896540
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp 1704896540
transform 1 0 4508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1704896540
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp 1704896540
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_61
timestamp 1704896540
transform 1 0 6164 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_73
timestamp 1704896540
transform 1 0 7268 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_79
timestamp 1704896540
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp 1704896540
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_85
timestamp 1704896540
transform 1 0 8372 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_93
timestamp 1704896540
transform 1 0 9108 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_97
timestamp 1704896540
transform 1 0 9476 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1704896540
transform 1 0 10580 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_116
timestamp 1704896540
transform 1 0 11224 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_128
timestamp 1704896540
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_133
timestamp 1704896540
transform 1 0 12788 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp 1704896540
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_141
timestamp 1704896540
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_147
timestamp 1704896540
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp 1704896540
transform 1 0 14444 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1704896540
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1704896540
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_172
timestamp 1704896540
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_187
timestamp 1704896540
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp 1704896540
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp 1704896540
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1704896540
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 3588 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 12328 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 2668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform 1 0 920 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 6532 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 6532 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 12328 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform 1 0 1932 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 4416 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform 1 0 12696 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16376 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform -1 0 14444 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform -1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1704896540
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 9200 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform -1 0 7820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1704896540
transform 1 0 2576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1704896540
transform 1 0 920 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1704896540
transform 1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp 1704896540
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp 1704896540
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp 1704896540
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp 1704896540
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp 1704896540
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1704896540
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp 1704896540
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1704896540
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp 1704896540
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1704896540
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 1704896540
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp 1704896540
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 1704896540
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 1704896540
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 1704896540
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 1704896540
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 1704896540
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 1704896540
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp 1704896540
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp 1704896540
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp 1704896540
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp 1704896540
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp 1704896540
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp 1704896540
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp 1704896540
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp 1704896540
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp 1704896540
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp 1704896540
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp 1704896540
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp 1704896540
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp 1704896540
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp 1704896540
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp 1704896540
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp 1704896540
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp 1704896540
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp 1704896540
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp 1704896540
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp 1704896540
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp 1704896540
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp 1704896540
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp 1704896540
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp 1704896540
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp 1704896540
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp 1704896540
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp 1704896540
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp 1704896540
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp 1704896540
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp 1704896540
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp 1704896540
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp 1704896540
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp 1704896540
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp 1704896540
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp 1704896540
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp 1704896540
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp 1704896540
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp 1704896540
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp 1704896540
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp 1704896540
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp 1704896540
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp 1704896540
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp 1704896540
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp 1704896540
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp 1704896540
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp 1704896540
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp 1704896540
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp 1704896540
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
<< labels >>
rlabel metal2 s 10061 19040 10061 19040 4 VGND
rlabel metal1 s 9982 18496 9982 18496 4 VPWR
rlabel metal2 s 16974 17918 16974 17918 4 _000_
rlabel metal2 s 4549 11186 4549 11186 4 _001_
rlabel metal2 s 6026 11458 6026 11458 4 _002_
rlabel metal2 s 4462 13634 4462 13634 4 _003_
rlabel metal2 s 6665 13838 6665 13838 4 _004_
rlabel metal1 s 4554 15674 4554 15674 4 _005_
rlabel metal1 s 4232 17306 4232 17306 4 _006_
rlabel metal1 s 2387 16694 2387 16694 4 _007_
rlabel metal1 s 1798 15538 1798 15538 4 _008_
rlabel metal1 s 2162 14042 2162 14042 4 _009_
rlabel metal2 s 1058 12988 1058 12988 4 _010_
rlabel metal1 s 3005 12682 3005 12682 4 _011_
rlabel metal2 s 4002 11492 4002 11492 4 _012_
rlabel metal1 s 8924 6698 8924 6698 4 _013_
rlabel metal2 s 9246 9180 9246 9180 4 _014_
rlabel metal1 s 9664 5746 9664 5746 4 _015_
rlabel metal1 s 9250 8398 9250 8398 4 _016_
rlabel metal1 s 9977 5134 9977 5134 4 _017_
rlabel metal1 s 11346 5814 11346 5814 4 _018_
rlabel metal2 s 11265 5066 11265 5066 4 _019_
rlabel metal2 s 11638 7480 11638 7480 4 _020_
rlabel metal2 s 11362 15844 11362 15844 4 _021_
rlabel metal2 s 15410 15164 15410 15164 4 _022_
rlabel metal1 s 13708 14586 13708 14586 4 _023_
rlabel metal2 s 15497 13838 15497 13838 4 _024_
rlabel metal1 s 11352 13838 11352 13838 4 _025_
rlabel metal1 s 10794 13430 10794 13430 4 _026_
rlabel metal2 s 14030 13158 14030 13158 4 _027_
rlabel metal1 s 11311 11662 11311 11662 4 _028_
rlabel metal1 s 18073 12750 18073 12750 4 _029_
rlabel metal1 s 8740 13158 8740 13158 4 _030_
rlabel metal1 s 8827 12682 8827 12682 4 _031_
rlabel metal2 s 9522 14722 9522 14722 4 _032_
rlabel metal2 s 10166 17408 10166 17408 4 _033_
rlabel metal2 s 9246 15810 9246 15810 4 _034_
rlabel metal2 s 8878 17986 8878 17986 4 _035_
rlabel metal1 s 7590 17850 7590 17850 4 _036_
rlabel metal1 s 7038 17306 7038 17306 4 _037_
rlabel metal1 s 2714 11764 2714 11764 4 _038_
rlabel metal1 s 4416 11866 4416 11866 4 _039_
rlabel metal1 s 4922 12104 4922 12104 4 _040_
rlabel metal1 s 4048 14450 4048 14450 4 _041_
rlabel metal2 s 5842 11628 5842 11628 4 _042_
rlabel metal1 s 4738 14382 4738 14382 4 _043_
rlabel metal1 s 4738 14280 4738 14280 4 _044_
rlabel metal2 s 4646 13804 4646 13804 4 _045_
rlabel metal1 s 5658 14314 5658 14314 4 _046_
rlabel metal1 s 5888 14246 5888 14246 4 _047_
rlabel metal1 s 6440 14450 6440 14450 4 _048_
rlabel metal1 s 4830 16150 4830 16150 4 _049_
rlabel metal1 s 4554 15572 4554 15572 4 _050_
rlabel metal1 s 3128 16014 3128 16014 4 _051_
rlabel metal1 s 4278 17102 4278 17102 4 _052_
rlabel metal1 s 2116 17102 2116 17102 4 _053_
rlabel metal2 s 3726 16898 3726 16898 4 _054_
rlabel metal2 s 1702 15742 1702 15742 4 _055_
rlabel metal1 s 2392 15062 2392 15062 4 _056_
rlabel metal2 s 2438 15096 2438 15096 4 _057_
rlabel metal1 s 2208 13838 2208 13838 4 _058_
rlabel metal1 s 2024 13498 2024 13498 4 _059_
rlabel metal1 s 1104 13362 1104 13362 4 _060_
rlabel metal1 s 3174 13838 3174 13838 4 _061_
rlabel metal1 s 2714 13872 2714 13872 4 _062_
rlabel metal1 s 3358 11594 3358 11594 4 _063_
rlabel metal2 s 8970 8942 8970 8942 4 _064_
rlabel metal1 s 10810 10608 10810 10608 4 _065_
rlabel metal2 s 10994 10404 10994 10404 4 _066_
rlabel metal1 s 10166 9418 10166 9418 4 _067_
rlabel metal2 s 17526 13634 17526 13634 4 _068_
rlabel metal1 s 16652 12682 16652 12682 4 _069_
rlabel metal1 s 12788 12614 12788 12614 4 _070_
rlabel metal1 s 13570 11696 13570 11696 4 _071_
rlabel metal1 s 13340 11730 13340 11730 4 _072_
rlabel metal2 s 17250 6766 17250 6766 4 _073_
rlabel metal1 s 15134 11628 15134 11628 4 _074_
rlabel metal1 s 17979 11254 17979 11254 4 _075_
rlabel metal1 s 17250 13974 17250 13974 4 _076_
rlabel metal1 s 16882 14586 16882 14586 4 _077_
rlabel metal2 s 17434 10540 17434 10540 4 _078_
rlabel metal1 s 16054 8466 16054 8466 4 _079_
rlabel metal2 s 15502 7004 15502 7004 4 _080_
rlabel metal1 s 16330 10098 16330 10098 4 _081_
rlabel metal1 s 15042 10506 15042 10506 4 _082_
rlabel metal2 s 15870 6800 15870 6800 4 _083_
rlabel metal1 s 14306 10132 14306 10132 4 _084_
rlabel metal2 s 16514 8806 16514 8806 4 _085_
rlabel metal1 s 15962 8364 15962 8364 4 _086_
rlabel metal1 s 14858 9962 14858 9962 4 _087_
rlabel metal1 s 15640 6290 15640 6290 4 _088_
rlabel metal1 s 14904 6426 14904 6426 4 _089_
rlabel metal2 s 18078 10370 18078 10370 4 _090_
rlabel metal1 s 16008 8534 16008 8534 4 _091_
rlabel metal2 s 17526 7548 17526 7548 4 _092_
rlabel metal1 s 17710 7922 17710 7922 4 _093_
rlabel metal1 s 17756 7514 17756 7514 4 _094_
rlabel metal1 s 15226 6834 15226 6834 4 _095_
rlabel metal2 s 15410 7650 15410 7650 4 _096_
rlabel metal1 s 15088 6358 15088 6358 4 _097_
rlabel metal1 s 15134 6630 15134 6630 4 _098_
rlabel metal2 s 14490 6494 14490 6494 4 _099_
rlabel metal1 s 9062 6800 9062 6800 4 _100_
rlabel metal2 s 12558 15878 12558 15878 4 _101_
rlabel metal2 s 15134 13634 15134 13634 4 _102_
rlabel metal1 s 15272 9418 15272 9418 4 _103_
rlabel metal1 s 14214 10030 14214 10030 4 _104_
rlabel metal2 s 12558 9010 12558 9010 4 _105_
rlabel metal1 s 11914 8466 11914 8466 4 _106_
rlabel metal1 s 17250 8908 17250 8908 4 _107_
rlabel metal1 s 14168 11118 14168 11118 4 _108_
rlabel metal1 s 16238 9622 16238 9622 4 _109_
rlabel metal2 s 14766 8959 14766 8959 4 _110_
rlabel metal2 s 11822 8704 11822 8704 4 _111_
rlabel metal2 s 10810 8840 10810 8840 4 _112_
rlabel metal1 s 14628 9146 14628 9146 4 _113_
rlabel metal2 s 13110 9180 13110 9180 4 _114_
rlabel metal2 s 12926 9316 12926 9316 4 _115_
rlabel metal1 s 11408 9486 11408 9486 4 _116_
rlabel metal1 s 9798 9554 9798 9554 4 _117_
rlabel metal1 s 10304 9146 10304 9146 4 _118_
rlabel metal1 s 10212 9486 10212 9486 4 _119_
rlabel metal1 s 13570 14892 13570 14892 4 _120_
rlabel metal2 s 9338 8942 9338 8942 4 _121_
rlabel metal1 s 16836 6222 16836 6222 4 _122_
rlabel metal1 s 17158 6426 17158 6426 4 _123_
rlabel metal1 s 17158 6324 17158 6324 4 _124_
rlabel metal1 s 14858 6154 14858 6154 4 _125_
rlabel metal1 s 14812 8058 14812 8058 4 _126_
rlabel metal1 s 14214 8364 14214 8364 4 _127_
rlabel metal1 s 13938 9588 13938 9588 4 _128_
rlabel metal2 s 14214 7378 14214 7378 4 _129_
rlabel metal1 s 14076 10438 14076 10438 4 _130_
rlabel metal1 s 15778 10166 15778 10166 4 _131_
rlabel metal2 s 14030 9724 14030 9724 4 _132_
rlabel metal1 s 14214 7276 14214 7276 4 _133_
rlabel metal2 s 14030 6698 14030 6698 4 _134_
rlabel metal1 s 14122 6698 14122 6698 4 _135_
rlabel metal1 s 13708 6222 13708 6222 4 _136_
rlabel metal1 s 10350 6358 10350 6358 4 _137_
rlabel metal1 s 9568 6426 9568 6426 4 _138_
rlabel metal2 s 10258 15237 10258 15237 4 _139_
rlabel metal1 s 13846 8942 13846 8942 4 _140_
rlabel metal1 s 14030 9010 14030 9010 4 _141_
rlabel metal2 s 13662 9248 13662 9248 4 _142_
rlabel metal1 s 16790 8058 16790 8058 4 _143_
rlabel metal1 s 13754 9588 13754 9588 4 _144_
rlabel metal1 s 14858 12818 14858 12818 4 _145_
rlabel metal2 s 15318 10812 15318 10812 4 _146_
rlabel metal1 s 14582 10064 14582 10064 4 _147_
rlabel metal1 s 14076 9554 14076 9554 4 _148_
rlabel metal1 s 10902 9554 10902 9554 4 _149_
rlabel metal1 s 9154 9452 9154 9452 4 _150_
rlabel metal1 s 10120 8058 10120 8058 4 _151_
rlabel metal2 s 12650 8908 12650 8908 4 _152_
rlabel metal1 s 12650 7956 12650 7956 4 _153_
rlabel metal2 s 12834 7718 12834 7718 4 _154_
rlabel metal2 s 12190 8228 12190 8228 4 _155_
rlabel metal1 s 11822 7854 11822 7854 4 _156_
rlabel metal1 s 10534 7922 10534 7922 4 _157_
rlabel metal3 s 10649 16660 10649 16660 4 _158_
rlabel metal1 s 12558 6766 12558 6766 4 _159_
rlabel metal1 s 11822 6766 11822 6766 4 _160_
rlabel metal1 s 10902 6222 10902 6222 4 _161_
rlabel metal1 s 10672 6834 10672 6834 4 _162_
rlabel metal2 s 10534 7004 10534 7004 4 _163_
rlabel metal1 s 11546 15436 11546 15436 4 _164_
rlabel metal1 s 13018 15130 13018 15130 4 _165_
rlabel metal1 s 14076 15946 14076 15946 4 _166_
rlabel metal2 s 12834 15776 12834 15776 4 _167_
rlabel metal1 s 15226 15572 15226 15572 4 _168_
rlabel metal1 s 14030 14926 14030 14926 4 _169_
rlabel metal2 s 12750 13430 12750 13430 4 _170_
rlabel metal1 s 13708 14926 13708 14926 4 _171_
rlabel metal2 s 13570 14620 13570 14620 4 _172_
rlabel metal1 s 15226 14450 15226 14450 4 _173_
rlabel metal2 s 11454 14178 11454 14178 4 _174_
rlabel metal1 s 13018 13260 13018 13260 4 _175_
rlabel metal2 s 13570 13022 13570 13022 4 _176_
rlabel metal2 s 10534 13158 10534 13158 4 _177_
rlabel metal1 s 14076 11866 14076 11866 4 _178_
rlabel metal1 s 11960 12750 11960 12750 4 _179_
rlabel metal1 s 11546 12614 11546 12614 4 _180_
rlabel metal2 s 17158 14620 17158 14620 4 _181_
rlabel metal1 s 14996 12886 14996 12886 4 _182_
rlabel metal2 s 18170 13872 18170 13872 4 _183_
rlabel metal1 s 9890 17204 9890 17204 4 _184_
rlabel metal2 s 8234 13124 8234 13124 4 _185_
rlabel metal1 s 9568 12410 9568 12410 4 _186_
rlabel metal1 s 8970 14586 8970 14586 4 _187_
rlabel metal1 s 9430 17170 9430 17170 4 _188_
rlabel metal1 s 9798 15674 9798 15674 4 _189_
rlabel metal1 s 8188 17850 8188 17850 4 _190_
rlabel metal1 s 6992 17850 6992 17850 4 _191_
rlabel metal1 s 7452 17170 7452 17170 4 _192_
rlabel metal1 s 9154 17544 9154 17544 4 _193_
rlabel metal2 s 7958 17408 7958 17408 4 _194_
rlabel metal1 s 8280 15334 8280 15334 4 _195_
rlabel metal1 s 6578 17238 6578 17238 4 _196_
rlabel metal1 s 7314 15674 7314 15674 4 _197_
rlabel metal2 s 12374 15674 12374 15674 4 _198_
rlabel metal1 s 7958 15436 7958 15436 4 _199_
rlabel metal1 s 7222 14586 7222 14586 4 _200_
rlabel metal1 s 7038 15912 7038 15912 4 _201_
rlabel metal1 s 6946 14450 6946 14450 4 _202_
rlabel metal1 s 7820 14586 7820 14586 4 _203_
rlabel metal2 s 7038 12070 7038 12070 4 _204_
rlabel metal1 s 6900 13158 6900 13158 4 _205_
rlabel metal1 s 6578 16082 6578 16082 4 _206_
rlabel metal2 s 7268 12580 7268 12580 4 _207_
rlabel metal2 s 7452 15436 7452 15436 4 _208_
rlabel metal1 s 7301 15538 7301 15538 4 _209_
rlabel metal2 s 13294 15742 13294 15742 4 _210_
rlabel metal1 s 12742 15572 12742 15572 4 _211_
rlabel metal2 s 6210 14824 6210 14824 4 _212_
rlabel metal3 s 18515 15980 18515 15980 4 clk
rlabel metal2 s 7130 13804 7130 13804 4 clknet_0_clk
rlabel metal2 s 2254 11764 2254 11764 4 clknet_2_0__leaf_clk
rlabel metal1 s 2208 15538 2208 15538 4 clknet_2_1__leaf_clk
rlabel metal2 s 9890 8670 9890 8670 4 clknet_2_2__leaf_clk
rlabel metal1 s 15226 14994 15226 14994 4 clknet_2_3__leaf_clk
rlabel metal1 s 18538 12954 18538 12954 4 cnt_zero
rlabel metal1 s 16054 18802 16054 18802 4 data[0]
rlabel metal1 s 14260 18802 14260 18802 4 data[1]
rlabel metal1 s 12604 18802 12604 18802 4 data[2]
rlabel metal1 s 11132 18802 11132 18802 4 data[3]
rlabel metal1 s 9200 18802 9200 18802 4 data[4]
rlabel metal1 s 7544 18802 7544 18802 4 data[5]
rlabel metal1 s 5888 18802 5888 18802 4 data[6]
rlabel metal1 s 4232 18802 4232 18802 4 data[7]
rlabel metal1 s 2576 18802 2576 18802 4 ext_data
rlabel metal1 s 920 18802 920 18802 4 load_divider
rlabel metal1 s 17572 18802 17572 18802 4 n_rst
rlabel metal1 s 12926 13362 12926 13362 4 net1
rlabel metal1 s 6992 17714 6992 17714 4 net10
rlabel metal1 s 17296 18190 17296 18190 4 net11
rlabel metal1 s 16146 17782 16146 17782 4 net12
rlabel metal1 s 3450 11662 3450 11662 4 net13
rlabel metal1 s 2622 13804 2622 13804 4 net14
rlabel metal1 s 11454 12206 11454 12206 4 net15
rlabel metal1 s 1426 13396 1426 13396 4 net16
rlabel metal1 s 1798 12342 1798 12342 4 net17
rlabel metal1 s 4462 15504 4462 15504 4 net18
rlabel metal1 s 5290 17102 5290 17102 4 net19
rlabel metal1 s 13018 12886 13018 12886 4 net2
rlabel metal1 s 11224 13362 11224 13362 4 net20
rlabel metal2 s 2622 15708 2622 15708 4 net21
rlabel metal1 s 3864 16218 3864 16218 4 net22
rlabel metal1 s 13478 13838 13478 13838 4 net23
rlabel metal2 s 12650 16558 12650 16558 4 net3
rlabel metal2 s 10258 18394 10258 18394 4 net4
rlabel metal2 s 9430 17068 9430 17068 4 net5
rlabel metal2 s 8694 18156 8694 18156 4 net6
rlabel metal2 s 7498 17578 7498 17578 4 net7
rlabel metal1 s 7314 17102 7314 17102 4 net8
rlabel metal1 s 9154 11220 9154 11220 4 net9
rlabel metal2 s 1242 1996 1242 1996 4 r2r_out[0]
rlabel metal1 s 5842 4114 5842 4114 4 r2r_out[1]
rlabel metal1 s 7452 3706 7452 3706 4 r2r_out[2]
rlabel metal2 s 8694 1557 8694 1557 4 r2r_out[3]
rlabel metal2 s 11178 1435 11178 1435 4 r2r_out[4]
rlabel metal1 s 13202 5542 13202 5542 4 r2r_out[5]
rlabel metal2 s 16146 2676 16146 2676 4 r2r_out[6]
rlabel metal1 s 18354 4998 18354 4998 4 r2r_out[7]
rlabel metal1 s 6394 13362 6394 13362 4 sine_lookup.count\[0\]
rlabel metal2 s 2622 12682 2622 12682 4 sine_lookup.count\[10\]
rlabel metal1 s 3358 11322 3358 11322 4 sine_lookup.count\[11\]
rlabel metal1 s 5520 12274 5520 12274 4 sine_lookup.count\[1\]
rlabel metal2 s 6762 14994 6762 14994 4 sine_lookup.count\[2\]
rlabel metal1 s 5520 14450 5520 14450 4 sine_lookup.count\[3\]
rlabel metal1 s 5566 16524 5566 16524 4 sine_lookup.count\[4\]
rlabel metal1 s 7406 15946 7406 15946 4 sine_lookup.count\[5\]
rlabel metal1 s 6762 15946 6762 15946 4 sine_lookup.count\[6\]
rlabel metal1 s 1794 16048 1794 16048 4 sine_lookup.count\[7\]
rlabel metal1 s 3450 14246 3450 14246 4 sine_lookup.count\[8\]
rlabel metal1 s 2438 12376 2438 12376 4 sine_lookup.count\[9\]
rlabel metal1 s 7498 12750 7498 12750 4 sine_lookup.divider\[0\]
rlabel metal1 s 9798 12614 9798 12614 4 sine_lookup.divider\[1\]
rlabel metal2 s 8142 14620 8142 14620 4 sine_lookup.divider\[2\]
rlabel metal1 s 10902 17714 10902 17714 4 sine_lookup.divider\[3\]
rlabel metal2 s 10074 16422 10074 16422 4 sine_lookup.divider\[4\]
rlabel metal1 s 9292 17102 9292 17102 4 sine_lookup.divider\[5\]
rlabel metal2 s 6302 17578 6302 17578 4 sine_lookup.divider\[6\]
rlabel metal1 s 6026 17136 6026 17136 4 sine_lookup.divider\[7\]
rlabel metal2 s 17894 17272 17894 17272 4 sine_lookup.rst
rlabel metal1 s 17296 14246 17296 14246 4 sine_lookup.sine_input\[0\]
rlabel metal1 s 17342 14450 17342 14450 4 sine_lookup.sine_input\[1\]
rlabel metal1 s 17013 13838 17013 13838 4 sine_lookup.sine_input\[2\]
rlabel metal2 s 16606 14246 16606 14246 4 sine_lookup.sine_input\[3\]
rlabel metal1 s 12650 12716 12650 12716 4 sine_lookup.sine_input\[4\]
rlabel metal1 s 12926 12852 12926 12852 4 sine_lookup.sine_input\[5\]
rlabel metal1 s 15410 13362 15410 13362 4 sine_lookup.sine_input\[6\]
rlabel metal2 s 10626 10353 10626 10353 4 sine_lookup.sine_input\[7\]
flabel metal4 s 19251 496 19571 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14536 496 14856 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9821 496 10141 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5106 496 5426 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16894 496 17214 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12179 496 12499 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7464 496 7784 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2749 496 3069 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 19062 19600 19118 20000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal3 s 19600 9800 20000 9920 0 FreeSans 600 0 0 0 cnt_zero
port 4 nsew
flabel metal2 s 15750 19600 15806 20000 0 FreeSans 280 90 0 0 data[0]
port 5 nsew
flabel metal2 s 14094 19600 14150 20000 0 FreeSans 280 90 0 0 data[1]
port 6 nsew
flabel metal2 s 12438 19600 12494 20000 0 FreeSans 280 90 0 0 data[2]
port 7 nsew
flabel metal2 s 10782 19600 10838 20000 0 FreeSans 280 90 0 0 data[3]
port 8 nsew
flabel metal2 s 9126 19600 9182 20000 0 FreeSans 280 90 0 0 data[4]
port 9 nsew
flabel metal2 s 7470 19600 7526 20000 0 FreeSans 280 90 0 0 data[5]
port 10 nsew
flabel metal2 s 5814 19600 5870 20000 0 FreeSans 280 90 0 0 data[6]
port 11 nsew
flabel metal2 s 4158 19600 4214 20000 0 FreeSans 280 90 0 0 data[7]
port 12 nsew
flabel metal2 s 2502 19600 2558 20000 0 FreeSans 280 90 0 0 ext_data
port 13 nsew
flabel metal2 s 846 19600 902 20000 0 FreeSans 280 90 0 0 load_divider
port 14 nsew
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 280 90 0 0 n_rst
port 15 nsew
flabel metal2 s 1214 0 1270 400 0 FreeSans 280 90 0 0 r2r_out[0]
port 16 nsew
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 r2r_out[1]
port 17 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 r2r_out[2]
port 18 nsew
flabel metal2 s 8666 0 8722 400 0 FreeSans 280 90 0 0 r2r_out[3]
port 19 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 r2r_out[4]
port 20 nsew
flabel metal2 s 13634 0 13690 400 0 FreeSans 280 90 0 0 r2r_out[5]
port 21 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 r2r_out[6]
port 22 nsew
flabel metal2 s 18602 0 18658 400 0 FreeSans 280 90 0 0 r2r_out[7]
port 23 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string GDS_END 1220090
string GDS_FILE ../gds/r2r_dac_control.gds
string GDS_START 443832
<< end >>
