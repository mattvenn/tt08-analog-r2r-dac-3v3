magic
tech sky130A
magscale 1 2
timestamp 1720527363
<< psubdiff >>
rect -1000 10700 -700 10724
rect -624 10700 -600 11100
rect 12900 10700 12924 11100
rect 13000 10700 13300 10724
rect -1000 976 -700 1000
rect 13000 976 13300 1000
<< psubdiffcont >>
rect -600 10700 12900 11100
rect -1000 1000 -700 10700
rect 13000 1000 13300 10700
<< locali >>
rect -1000 10700 -700 10716
rect -616 10700 -600 11100
rect 12900 10700 12916 11100
rect 13000 10700 13300 10716
rect -1000 984 -700 1000
rect 13000 984 13300 1000
<< viali >>
rect -500 10800 12800 11000
rect -900 1200 -800 10500
rect 13100 1200 13200 10500
<< metal1 >>
rect -1000 11000 13300 11100
rect -1000 10800 -500 11000
rect 12800 10800 13300 11000
rect -1000 10700 13300 10800
rect -1000 10500 -600 10700
rect -1000 1800 -900 10500
rect -800 10400 -600 10500
rect 12900 10500 13300 10700
rect 12900 10400 13100 10500
rect -800 10000 -200 10400
rect 0 10000 800 10400
rect 1000 10000 1800 10400
rect -800 1800 -700 10000
rect 2000 5700 2300 10400
rect 2500 10000 3300 10400
rect 3500 5700 3800 10400
rect 4000 10000 4800 10400
rect 5000 5700 5300 10400
rect 5500 10000 6300 10400
rect 6500 5700 6800 10400
rect 7000 10000 7800 10400
rect 8000 5700 8300 10400
rect 8500 10000 9300 10400
rect 9500 5700 9800 10400
rect 10000 10000 10800 10400
rect 11000 5700 11300 10400
rect 11500 10000 12300 10400
rect 12500 10000 13100 10400
rect 1000 5400 2300 5700
rect 2500 5400 3800 5700
rect 4000 5400 5300 5700
rect 5500 5400 6800 5700
rect 7000 5400 8300 5700
rect 8500 5400 9800 5700
rect 10000 5400 11300 5700
rect -1010 1500 -1000 1800
rect -700 1500 -690 1800
rect -1000 1200 -900 1500
rect -800 1200 -700 1500
rect -1000 1000 -700 1200
rect 1000 1000 1300 5400
rect 1490 1500 1500 1800
rect 1800 1500 1810 1800
rect -1000 600 -200 1000
rect 0 300 300 1000
rect 500 600 1300 1000
rect 1500 300 1800 1500
rect 2500 1000 2800 5400
rect 4000 1000 4300 5400
rect 5500 1000 5800 5400
rect 7000 1000 7300 5400
rect 8500 1000 8800 5400
rect 10000 1000 10300 5400
rect 13000 1200 13100 10000
rect 13200 1200 13300 10500
rect 13000 1000 13300 1200
rect 2000 600 2800 1000
rect 3000 300 3300 1000
rect 3500 600 4300 1000
rect 4500 300 4800 1000
rect 5000 600 5800 1000
rect 6000 300 6300 1000
rect 6500 600 7300 1000
rect 7500 300 7800 1000
rect 8000 600 8800 1000
rect 9000 300 9300 1000
rect 9500 600 10300 1000
rect 10500 300 10800 1000
rect 11000 600 11800 1000
rect 11300 300 11600 600
rect 12000 300 12300 1000
rect 12500 600 13300 1000
<< via1 >>
rect -1000 1500 -900 1800
rect -900 1500 -800 1800
rect -800 1500 -700 1800
rect 1500 1500 1800 1800
<< metal2 >>
rect -1000 1800 -700 1810
rect 1500 1800 1800 1810
rect -700 1500 1500 1800
rect -1000 1490 -700 1500
rect 1500 1490 1800 1500
use sky130_fd_pr__res_high_po_1p41_BF4AJ4  sky130_fd_pr__res_high_po_1p41_BF4AJ4_0
array 0 24 500 0 0 10000
timestamp 1720520928
transform 1 0 141 0 1 5516
box -141 -4916 141 4916
use sky130_fd_pr__res_high_po_1p41_NAL9NH  sky130_fd_pr__res_high_po_1p41_NAL9NH_0
timestamp 1720521380
transform 1 0 12641 0 1 5516
box -141 -4916 141 4916
use sky130_fd_pr__res_high_po_1p41_NAL9NH  sky130_fd_pr__res_high_po_1p41_NAL9NH_1
timestamp 1720521380
transform 1 0 -359 0 1 5516
box -141 -4916 141 4916
<< labels >>
flabel metal1 1500 300 1700 500 0 FreeSans 256 0 0 0 VGND
port 9 nsew
flabel metal1 3000 300 3200 500 0 FreeSans 256 0 0 0 b1
port 2 nsew
flabel metal1 0 300 200 500 0 FreeSans 256 0 0 0 b0
port 3 nsew
flabel metal1 4500 300 4700 500 0 FreeSans 256 0 0 0 b2
port 1 nsew
flabel metal1 6000 300 6200 500 0 FreeSans 256 0 0 0 b3
port 7 nsew
flabel metal1 7500 300 7700 500 0 FreeSans 256 0 0 0 b4
port 0 nsew
flabel metal1 9000 300 9200 500 0 FreeSans 256 0 0 0 b5
port 4 nsew
flabel metal1 10500 300 10700 500 0 FreeSans 256 0 0 0 b6
port 5 nsew
flabel metal1 12000 300 12200 500 0 FreeSans 256 0 0 0 b7
port 6 nsew
flabel metal1 11300 300 11500 500 0 FreeSans 256 0 0 0 out
port 8 nsew
flabel metal1 500 600 1300 1000 0 FreeSans 1600 0 0 0 a
flabel metal1 2000 600 2800 1000 0 FreeSans 1600 0 0 0 b
flabel metal1 3500 600 4300 1000 0 FreeSans 1600 0 0 0 c
flabel metal1 5000 600 5800 1000 0 FreeSans 1600 0 0 0 d
flabel metal1 6500 600 7300 1000 0 FreeSans 1600 0 0 0 e
flabel metal1 8000 600 8800 1000 0 FreeSans 1600 0 0 0 f
flabel metal1 9500 600 10300 1000 0 FreeSans 1600 0 0 0 g
<< end >>
