magic
tech sky130A
magscale 1 2
timestamp 1720438358
<< viali >>
rect 4445 18921 4479 18955
rect 949 18785 983 18819
rect 2605 18785 2639 18819
rect 4261 18785 4295 18819
rect 5917 18785 5951 18819
rect 7573 18785 7607 18819
rect 9229 18785 9263 18819
rect 9413 18785 9447 18819
rect 9689 18785 9723 18819
rect 11161 18785 11195 18819
rect 12725 18785 12759 18819
rect 14381 18785 14415 18819
rect 16313 18785 16347 18819
rect 17693 18785 17727 18819
rect 1225 18717 1259 18751
rect 2789 18649 2823 18683
rect 7757 18649 7791 18683
rect 14197 18649 14231 18683
rect 6101 18581 6135 18615
rect 9321 18581 9355 18615
rect 9505 18581 9539 18615
rect 10977 18581 11011 18615
rect 12541 18581 12575 18615
rect 16129 18581 16163 18615
rect 17509 18581 17543 18615
rect 11437 18377 11471 18411
rect 6285 18241 6319 18275
rect 8217 18241 8251 18275
rect 9137 18241 9171 18275
rect 9873 18241 9907 18275
rect 3617 18173 3651 18207
rect 5825 18173 5859 18207
rect 6377 18173 6411 18207
rect 8769 18173 8803 18207
rect 8861 18173 8895 18207
rect 9505 18173 9539 18207
rect 9597 18173 9631 18207
rect 11345 18173 11379 18207
rect 16773 18173 16807 18207
rect 5580 18105 5614 18139
rect 6101 18105 6135 18139
rect 7972 18105 8006 18139
rect 9045 18105 9079 18139
rect 9781 18105 9815 18139
rect 10118 18105 10152 18139
rect 3433 18037 3467 18071
rect 4445 18037 4479 18071
rect 6745 18037 6779 18071
rect 6837 18037 6871 18071
rect 8401 18037 8435 18071
rect 11253 18037 11287 18071
rect 14933 18037 14967 18071
rect 16681 18037 16715 18071
rect 2973 17833 3007 17867
rect 6193 17833 6227 17867
rect 8493 17833 8527 17867
rect 9045 17833 9079 17867
rect 15945 17833 15979 17867
rect 14473 17765 14507 17799
rect 1860 17697 1894 17731
rect 3065 17697 3099 17731
rect 3332 17697 3366 17731
rect 5089 17697 5123 17731
rect 6745 17697 6779 17731
rect 7941 17697 7975 17731
rect 9413 17697 9447 17731
rect 9505 17697 9539 17731
rect 9689 17697 9723 17731
rect 10609 17697 10643 17731
rect 11621 17697 11655 17731
rect 1593 17629 1627 17663
rect 4997 17629 5031 17663
rect 6469 17629 6503 17663
rect 8217 17629 8251 17663
rect 9321 17629 9355 17663
rect 14197 17629 14231 17663
rect 4445 17493 4479 17527
rect 5457 17493 5491 17527
rect 6653 17493 6687 17527
rect 8309 17493 8343 17527
rect 9321 17493 9355 17527
rect 9597 17493 9631 17527
rect 10517 17493 10551 17527
rect 11437 17493 11471 17527
rect 2421 17289 2455 17323
rect 2697 17289 2731 17323
rect 3525 17289 3559 17323
rect 6561 17289 6595 17323
rect 10793 17289 10827 17323
rect 3893 17153 3927 17187
rect 4445 17153 4479 17187
rect 4721 17153 4755 17187
rect 1777 17085 1811 17119
rect 1961 17085 1995 17119
rect 2053 17085 2087 17119
rect 2237 17085 2271 17119
rect 3709 17085 3743 17119
rect 4353 17085 4387 17119
rect 4905 17085 4939 17119
rect 4998 17085 5032 17119
rect 5273 17085 5307 17119
rect 5411 17085 5445 17119
rect 5641 17085 5675 17119
rect 5789 17085 5823 17119
rect 6009 17085 6043 17119
rect 6125 17085 6159 17119
rect 6653 17085 6687 17119
rect 8125 17085 8159 17119
rect 9229 17085 9263 17119
rect 10701 17085 10735 17119
rect 2665 17017 2699 17051
rect 2881 17017 2915 17051
rect 5181 17017 5215 17051
rect 5917 17017 5951 17051
rect 7858 17017 7892 17051
rect 9496 17017 9530 17051
rect 1869 16949 1903 16983
rect 2513 16949 2547 16983
rect 5549 16949 5583 16983
rect 6285 16949 6319 16983
rect 6745 16949 6779 16983
rect 10609 16949 10643 16983
rect 2329 16745 2363 16779
rect 3985 16745 4019 16779
rect 7113 16745 7147 16779
rect 7205 16745 7239 16779
rect 7849 16745 7883 16779
rect 9045 16745 9079 16779
rect 9137 16745 9171 16779
rect 9781 16745 9815 16779
rect 12081 16745 12115 16779
rect 5825 16677 5859 16711
rect 9965 16677 9999 16711
rect 2513 16609 2547 16643
rect 4077 16609 4111 16643
rect 5181 16609 5215 16643
rect 5365 16609 5399 16643
rect 6009 16609 6043 16643
rect 6101 16609 6135 16643
rect 6377 16609 6411 16643
rect 6469 16609 6503 16643
rect 6745 16609 6779 16643
rect 6837 16609 6871 16643
rect 8309 16609 8343 16643
rect 8677 16609 8711 16643
rect 8861 16609 8895 16643
rect 9597 16609 9631 16643
rect 9873 16609 9907 16643
rect 10057 16609 10091 16643
rect 11161 16609 11195 16643
rect 11805 16609 11839 16643
rect 11897 16609 11931 16643
rect 12449 16609 12483 16643
rect 5273 16541 5307 16575
rect 5457 16541 5491 16575
rect 7573 16541 7607 16575
rect 7665 16541 7699 16575
rect 9505 16541 9539 16575
rect 11621 16541 11655 16575
rect 11713 16541 11747 16575
rect 12265 16541 12299 16575
rect 12357 16541 12391 16575
rect 12541 16541 12575 16575
rect 5641 16473 5675 16507
rect 6653 16473 6687 16507
rect 8493 16473 8527 16507
rect 11345 16473 11379 16507
rect 6285 16405 6319 16439
rect 6745 16405 6779 16439
rect 8861 16405 8895 16439
rect 11437 16405 11471 16439
rect 4813 16201 4847 16235
rect 8953 16201 8987 16235
rect 9413 16133 9447 16167
rect 9781 16133 9815 16167
rect 4537 16065 4571 16099
rect 7113 16065 7147 16099
rect 8769 16065 8803 16099
rect 10793 16065 10827 16099
rect 13553 16065 13587 16099
rect 1869 15997 1903 16031
rect 2053 15997 2087 16031
rect 2145 15997 2179 16031
rect 2697 15997 2731 16031
rect 4445 15997 4479 16031
rect 7021 15997 7055 16031
rect 9045 15997 9079 16031
rect 9413 15997 9447 16031
rect 9597 15997 9631 16031
rect 9689 15997 9723 16031
rect 10057 15997 10091 16031
rect 11161 15997 11195 16031
rect 11345 15997 11379 16031
rect 11621 15997 11655 16031
rect 11897 15997 11931 16031
rect 13829 15997 13863 16031
rect 2513 15929 2547 15963
rect 9781 15929 9815 15963
rect 11805 15929 11839 15963
rect 12142 15929 12176 15963
rect 1685 15861 1719 15895
rect 2881 15861 2915 15895
rect 6837 15861 6871 15895
rect 7481 15861 7515 15895
rect 8493 15861 8527 15895
rect 9965 15861 9999 15895
rect 10241 15861 10275 15895
rect 13277 15861 13311 15895
rect 15117 15861 15151 15895
rect 1133 15657 1167 15691
rect 1961 15657 1995 15691
rect 2421 15657 2455 15691
rect 10517 15657 10551 15691
rect 11345 15657 11379 15691
rect 13093 15657 13127 15691
rect 1317 15589 1351 15623
rect 1777 15589 1811 15623
rect 2053 15589 2087 15623
rect 9404 15589 9438 15623
rect 857 15521 891 15555
rect 2145 15521 2179 15555
rect 3534 15521 3568 15555
rect 3801 15521 3835 15555
rect 6929 15521 6963 15555
rect 8677 15521 8711 15555
rect 10793 15521 10827 15555
rect 11161 15521 11195 15555
rect 11437 15521 11471 15555
rect 11621 15521 11655 15555
rect 11805 15521 11839 15555
rect 11989 15521 12023 15555
rect 12265 15521 12299 15555
rect 12633 15521 12667 15555
rect 12909 15521 12943 15555
rect 1685 15453 1719 15487
rect 9137 15453 9171 15487
rect 10977 15453 11011 15487
rect 1041 15317 1075 15351
rect 1317 15317 1351 15351
rect 2329 15317 2363 15351
rect 10701 15317 10735 15351
rect 11437 15317 11471 15351
rect 11897 15317 11931 15351
rect 2881 15113 2915 15147
rect 3433 15113 3467 15147
rect 8401 15113 8435 15147
rect 11529 15113 11563 15147
rect 11713 15113 11747 15147
rect 3065 15045 3099 15079
rect 857 14977 891 15011
rect 1124 14909 1158 14943
rect 2513 14909 2547 14943
rect 3249 14909 3283 14943
rect 3617 14909 3651 14943
rect 3801 14909 3835 14943
rect 4077 14909 4111 14943
rect 4261 14909 4295 14943
rect 4905 14909 4939 14943
rect 6285 14909 6319 14943
rect 6552 14909 6586 14943
rect 9781 14909 9815 14943
rect 14841 14909 14875 14943
rect 14933 14909 14967 14943
rect 4445 14841 4479 14875
rect 4721 14841 4755 14875
rect 9514 14841 9548 14875
rect 11345 14841 11379 14875
rect 11561 14841 11595 14875
rect 2237 14773 2271 14807
rect 2881 14773 2915 14807
rect 3985 14773 4019 14807
rect 5089 14773 5123 14807
rect 7665 14773 7699 14807
rect 15485 14773 15519 14807
rect 3985 14569 4019 14603
rect 5825 14569 5859 14603
rect 7849 14569 7883 14603
rect 8309 14569 8343 14603
rect 8953 14569 8987 14603
rect 2129 14501 2163 14535
rect 2329 14501 2363 14535
rect 4169 14501 4203 14535
rect 5273 14501 5307 14535
rect 4537 14433 4571 14467
rect 4813 14433 4847 14467
rect 6938 14433 6972 14467
rect 7205 14433 7239 14467
rect 7297 14433 7331 14467
rect 8769 14433 8803 14467
rect 11621 14433 11655 14467
rect 11989 14433 12023 14467
rect 12173 14433 12207 14467
rect 12265 14433 12299 14467
rect 12449 14433 12483 14467
rect 12716 14433 12750 14467
rect 14933 14433 14967 14467
rect 15209 14433 15243 14467
rect 7573 14365 7607 14399
rect 8677 14365 8711 14399
rect 11897 14365 11931 14399
rect 1961 14297 1995 14331
rect 4905 14297 4939 14331
rect 11713 14297 11747 14331
rect 2145 14229 2179 14263
rect 4169 14229 4203 14263
rect 4629 14229 4663 14263
rect 5273 14229 5307 14263
rect 5457 14229 5491 14263
rect 7665 14229 7699 14263
rect 11621 14229 11655 14263
rect 11989 14229 12023 14263
rect 13829 14229 13863 14263
rect 3341 14025 3375 14059
rect 4997 14025 5031 14059
rect 5549 14025 5583 14059
rect 11253 14025 11287 14059
rect 12081 14025 12115 14059
rect 12541 14025 12575 14059
rect 12909 14025 12943 14059
rect 11437 13957 11471 13991
rect 13921 13957 13955 13991
rect 4721 13889 4755 13923
rect 6653 13889 6687 13923
rect 6929 13889 6963 13923
rect 12449 13889 12483 13923
rect 1685 13821 1719 13855
rect 1869 13821 1903 13855
rect 2053 13821 2087 13855
rect 2145 13821 2179 13855
rect 2973 13821 3007 13855
rect 4465 13821 4499 13855
rect 5365 13821 5399 13855
rect 6561 13821 6595 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 10885 13821 10919 13855
rect 11161 13821 11195 13855
rect 11897 13821 11931 13855
rect 12173 13821 12207 13855
rect 12725 13821 12759 13855
rect 14013 13821 14047 13855
rect 16221 13821 16255 13855
rect 16497 13821 16531 13855
rect 4813 13753 4847 13787
rect 11069 13753 11103 13787
rect 11437 13753 11471 13787
rect 2329 13685 2363 13719
rect 5013 13685 5047 13719
rect 5181 13685 5215 13719
rect 9965 13685 9999 13719
rect 10701 13685 10735 13719
rect 11713 13685 11747 13719
rect 2605 13481 2639 13515
rect 7757 13481 7791 13515
rect 11713 13481 11747 13515
rect 1308 13413 1342 13447
rect 4997 13413 5031 13447
rect 5181 13413 5215 13447
rect 8585 13413 8619 13447
rect 8769 13413 8803 13447
rect 12326 13413 12360 13447
rect 2513 13345 2547 13379
rect 2789 13345 2823 13379
rect 2973 13345 3007 13379
rect 6009 13345 6043 13379
rect 7481 13345 7515 13379
rect 8033 13345 8067 13379
rect 8401 13345 8435 13379
rect 9321 13345 9355 13379
rect 9588 13345 9622 13379
rect 11713 13345 11747 13379
rect 11805 13345 11839 13379
rect 11989 13345 12023 13379
rect 14933 13345 14967 13379
rect 15117 13345 15151 13379
rect 16221 13345 16255 13379
rect 16589 13345 16623 13379
rect 1041 13277 1075 13311
rect 5825 13277 5859 13311
rect 7665 13277 7699 13311
rect 8309 13277 8343 13311
rect 11529 13277 11563 13311
rect 12081 13277 12115 13311
rect 10701 13209 10735 13243
rect 15301 13209 15335 13243
rect 2421 13141 2455 13175
rect 6193 13141 6227 13175
rect 10977 13141 11011 13175
rect 13461 13141 13495 13175
rect 17877 13141 17911 13175
rect 3985 12937 4019 12971
rect 4445 12937 4479 12971
rect 5641 12937 5675 12971
rect 8033 12937 8067 12971
rect 9965 12937 9999 12971
rect 10333 12937 10367 12971
rect 11253 12937 11287 12971
rect 12817 12937 12851 12971
rect 9505 12869 9539 12903
rect 10793 12869 10827 12903
rect 10425 12801 10459 12835
rect 1225 12733 1259 12767
rect 2697 12733 2731 12767
rect 2881 12733 2915 12767
rect 3801 12733 3835 12767
rect 4169 12733 4203 12767
rect 4261 12733 4295 12767
rect 4905 12733 4939 12767
rect 6929 12733 6963 12767
rect 7205 12733 7239 12767
rect 7941 12733 7975 12767
rect 8125 12733 8159 12767
rect 8401 12733 8435 12767
rect 9505 12733 9539 12767
rect 9781 12733 9815 12767
rect 10149 12733 10183 12767
rect 10517 12733 10551 12767
rect 11069 12733 11103 12767
rect 11345 12733 11379 12767
rect 14197 12733 14231 12767
rect 14841 12733 14875 12767
rect 15117 12733 15151 12767
rect 1492 12665 1526 12699
rect 2789 12665 2823 12699
rect 3985 12665 4019 12699
rect 4721 12665 4755 12699
rect 10793 12665 10827 12699
rect 11529 12665 11563 12699
rect 13645 12665 13679 12699
rect 2605 12597 2639 12631
rect 3249 12597 3283 12631
rect 5089 12597 5123 12631
rect 7021 12597 7055 12631
rect 8585 12597 8619 12631
rect 9689 12597 9723 12631
rect 10609 12597 10643 12631
rect 10885 12597 10919 12631
rect 2421 12393 2455 12427
rect 2584 12393 2618 12427
rect 2881 12393 2915 12427
rect 5457 12393 5491 12427
rect 5825 12393 5859 12427
rect 12725 12393 12759 12427
rect 2789 12325 2823 12359
rect 14013 12325 14047 12359
rect 14933 12325 14967 12359
rect 3157 12257 3191 12291
rect 4169 12257 4203 12291
rect 4629 12257 4663 12291
rect 4813 12257 4847 12291
rect 6949 12257 6983 12291
rect 7205 12257 7239 12291
rect 7757 12257 7791 12291
rect 10333 12257 10367 12291
rect 10425 12257 10459 12291
rect 10977 12257 11011 12291
rect 11233 12257 11267 12291
rect 12817 12257 12851 12291
rect 13369 12257 13403 12291
rect 13645 12257 13679 12291
rect 14105 12257 14139 12291
rect 2881 12189 2915 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 5089 12189 5123 12223
rect 8033 12189 8067 12223
rect 9321 12189 9355 12223
rect 10057 12189 10091 12223
rect 10517 12189 10551 12223
rect 10609 12189 10643 12223
rect 5641 12121 5675 12155
rect 12357 12121 12391 12155
rect 2605 12053 2639 12087
rect 3065 12053 3099 12087
rect 3985 12053 4019 12087
rect 4445 12053 4479 12087
rect 5457 12053 5491 12087
rect 9505 12053 9539 12087
rect 10793 12053 10827 12087
rect 2697 11849 2731 11883
rect 4905 11849 4939 11883
rect 5181 11849 5215 11883
rect 5457 11849 5491 11883
rect 7665 11849 7699 11883
rect 10885 11849 10919 11883
rect 16221 11849 16255 11883
rect 2329 11713 2363 11747
rect 6285 11713 6319 11747
rect 2513 11645 2547 11679
rect 3525 11645 3559 11679
rect 5917 11645 5951 11679
rect 6101 11645 6135 11679
rect 10609 11645 10643 11679
rect 10701 11645 10735 11679
rect 10885 11645 10919 11679
rect 13645 11645 13679 11679
rect 15209 11645 15243 11679
rect 15393 11645 15427 11679
rect 16129 11645 16163 11679
rect 16405 11645 16439 11679
rect 3792 11577 3826 11611
rect 4997 11577 5031 11611
rect 5213 11577 5247 11611
rect 5641 11577 5675 11611
rect 5825 11577 5859 11611
rect 6552 11577 6586 11611
rect 14381 11577 14415 11611
rect 5365 11509 5399 11543
rect 5917 11509 5951 11543
rect 9321 11509 9355 11543
rect 15301 11509 15335 11543
rect 16681 11509 16715 11543
rect 2145 11305 2179 11339
rect 4077 11305 4111 11339
rect 4261 11305 4295 11339
rect 4705 11305 4739 11339
rect 6653 11305 6687 11339
rect 8217 11305 8251 11339
rect 8493 11305 8527 11339
rect 10057 11305 10091 11339
rect 10215 11305 10249 11339
rect 15853 11305 15887 11339
rect 2329 11237 2363 11271
rect 2789 11237 2823 11271
rect 4905 11237 4939 11271
rect 8309 11237 8343 11271
rect 10425 11237 10459 11271
rect 2053 11169 2087 11203
rect 2697 11169 2731 11203
rect 2973 11169 3007 11203
rect 3157 11169 3191 11203
rect 3709 11169 3743 11203
rect 6469 11169 6503 11203
rect 8401 11169 8435 11203
rect 8677 11169 8711 11203
rect 8861 11169 8895 11203
rect 8953 11169 8987 11203
rect 9229 11169 9263 11203
rect 9689 11169 9723 11203
rect 9781 11169 9815 11203
rect 11897 11169 11931 11203
rect 12633 11169 12667 11203
rect 14013 11169 14047 11203
rect 14197 11169 14231 11203
rect 14657 11169 14691 11203
rect 14749 11169 14783 11203
rect 14841 11169 14875 11203
rect 14959 11169 14993 11203
rect 15117 11169 15151 11203
rect 15485 11169 15519 11203
rect 15669 11169 15703 11203
rect 15761 11169 15795 11203
rect 15945 11169 15979 11203
rect 16313 11169 16347 11203
rect 16405 11169 16439 11203
rect 16589 11169 16623 11203
rect 16773 11169 16807 11203
rect 16865 11169 16899 11203
rect 16957 11169 16991 11203
rect 17141 11169 17175 11203
rect 8033 11101 8067 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 15577 11101 15611 11135
rect 4537 11033 4571 11067
rect 8309 11033 8343 11067
rect 9965 11033 9999 11067
rect 14013 11033 14047 11067
rect 16129 11033 16163 11067
rect 16497 11033 16531 11067
rect 17141 11033 17175 11067
rect 1869 10965 1903 10999
rect 2329 10965 2363 10999
rect 4077 10965 4111 10999
rect 4721 10965 4755 10999
rect 9045 10965 9079 10999
rect 10241 10965 10275 10999
rect 14473 10965 14507 10999
rect 3065 10761 3099 10795
rect 9781 10761 9815 10795
rect 14105 10761 14139 10795
rect 14473 10761 14507 10795
rect 11805 10693 11839 10727
rect 17141 10693 17175 10727
rect 11345 10625 11379 10659
rect 16497 10625 16531 10659
rect 16589 10625 16623 10659
rect 1685 10557 1719 10591
rect 1952 10557 1986 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 8401 10557 8435 10591
rect 8668 10557 8702 10591
rect 11437 10557 11471 10591
rect 13553 10557 13587 10591
rect 13737 10557 13771 10591
rect 13829 10557 13863 10591
rect 14013 10567 14047 10601
rect 14289 10557 14323 10591
rect 14565 10557 14599 10591
rect 14841 10557 14875 10591
rect 14933 10557 14967 10591
rect 15025 10557 15059 10591
rect 15117 10557 15151 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 16957 10557 16991 10591
rect 7757 10421 7791 10455
rect 13553 10421 13587 10455
rect 13921 10421 13955 10455
rect 14657 10421 14691 10455
rect 15853 10421 15887 10455
rect 16037 10421 16071 10455
rect 16405 10421 16439 10455
rect 7021 10217 7055 10251
rect 14197 10217 14231 10251
rect 14289 10217 14323 10251
rect 17785 10217 17819 10251
rect 17877 10217 17911 10251
rect 10425 10149 10459 10183
rect 14565 10149 14599 10183
rect 16129 10149 16163 10183
rect 6929 10081 6963 10115
rect 7113 10081 7147 10115
rect 7389 10081 7423 10115
rect 7573 10081 7607 10115
rect 9873 10081 9907 10115
rect 10057 10081 10091 10115
rect 10241 10081 10275 10115
rect 11253 10081 11287 10115
rect 11989 10081 12023 10115
rect 13185 10081 13219 10115
rect 13277 10081 13311 10115
rect 13369 10081 13403 10115
rect 13645 10081 13679 10115
rect 14473 10081 14507 10115
rect 14749 10081 14783 10115
rect 16313 10081 16347 10115
rect 16405 10081 16439 10115
rect 9781 10013 9815 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 13921 10013 13955 10047
rect 14013 10013 14047 10047
rect 14381 10013 14415 10047
rect 17969 10013 18003 10047
rect 12909 9945 12943 9979
rect 14749 9945 14783 9979
rect 7481 9877 7515 9911
rect 10517 9877 10551 9911
rect 13001 9877 13035 9911
rect 16129 9877 16163 9911
rect 17417 9877 17451 9911
rect 10517 9673 10551 9707
rect 13829 9673 13863 9707
rect 14105 9673 14139 9707
rect 7941 9537 7975 9571
rect 9137 9537 9171 9571
rect 10333 9537 10367 9571
rect 11069 9537 11103 9571
rect 11897 9537 11931 9571
rect 8953 9469 8987 9503
rect 9689 9469 9723 9503
rect 9873 9469 9907 9503
rect 9965 9469 9999 9503
rect 10057 9469 10091 9503
rect 10417 9469 10451 9503
rect 13737 9469 13771 9503
rect 13921 9469 13955 9503
rect 14013 9469 14047 9503
rect 14197 9469 14231 9503
rect 15945 9469 15979 9503
rect 16037 9469 16071 9503
rect 16313 9469 16347 9503
rect 16405 9469 16439 9503
rect 7674 9401 7708 9435
rect 16129 9401 16163 9435
rect 6561 9333 6595 9367
rect 8493 9333 8527 9367
rect 8861 9333 8895 9367
rect 13553 9333 13587 9367
rect 15761 9333 15795 9367
rect 7481 9129 7515 9163
rect 9045 9129 9079 9163
rect 10241 9129 10275 9163
rect 13277 9129 13311 9163
rect 15853 9129 15887 9163
rect 16129 9129 16163 9163
rect 16957 9129 16991 9163
rect 17325 9129 17359 9163
rect 7665 9061 7699 9095
rect 8861 9061 8895 9095
rect 11989 9061 12023 9095
rect 12449 9061 12483 9095
rect 17969 9061 18003 9095
rect 7389 8993 7423 9027
rect 9137 8993 9171 9027
rect 9505 8993 9539 9027
rect 9689 8993 9723 9027
rect 9965 8993 9999 9027
rect 10333 8993 10367 9027
rect 10517 8993 10551 9027
rect 11621 8993 11655 9027
rect 11805 8993 11839 9027
rect 11897 8993 11931 9027
rect 12265 8993 12299 9027
rect 13093 8993 13127 9027
rect 13185 8993 13219 9027
rect 13553 8993 13587 9027
rect 15669 8993 15703 9027
rect 15945 8993 15979 9027
rect 16681 8993 16715 9027
rect 18153 8993 18187 9027
rect 9321 8925 9355 8959
rect 9781 8925 9815 8959
rect 12081 8925 12115 8959
rect 13461 8925 13495 8959
rect 16405 8925 16439 8959
rect 17417 8925 17451 8959
rect 17601 8925 17635 8959
rect 17785 8925 17819 8959
rect 7665 8857 7699 8891
rect 9597 8857 9631 8891
rect 11621 8857 11655 8891
rect 8861 8789 8895 8823
rect 10057 8789 10091 8823
rect 12173 8789 12207 8823
rect 12817 8789 12851 8823
rect 15669 8789 15703 8823
rect 16313 8789 16347 8823
rect 12265 8585 12299 8619
rect 13277 8585 13311 8619
rect 16313 8585 16347 8619
rect 17417 8585 17451 8619
rect 18337 8585 18371 8619
rect 8493 8517 8527 8551
rect 17509 8517 17543 8551
rect 13737 8449 13771 8483
rect 15209 8449 15243 8483
rect 15393 8449 15427 8483
rect 18061 8449 18095 8483
rect 9873 8381 9907 8415
rect 11989 8381 12023 8415
rect 12449 8381 12483 8415
rect 12725 8381 12759 8415
rect 13185 8381 13219 8415
rect 13369 8381 13403 8415
rect 13921 8381 13955 8415
rect 14197 8381 14231 8415
rect 14473 8381 14507 8415
rect 14657 8381 14691 8415
rect 14749 8381 14783 8415
rect 15117 8381 15151 8415
rect 15301 8381 15335 8415
rect 15761 8381 15795 8415
rect 15853 8381 15887 8415
rect 16037 8381 16071 8415
rect 16129 8381 16163 8415
rect 16497 8381 16531 8415
rect 16773 8381 16807 8415
rect 16921 8381 16955 8415
rect 17141 8381 17175 8415
rect 17279 8381 17313 8415
rect 17877 8381 17911 8415
rect 18337 8381 18371 8415
rect 18521 8381 18555 8415
rect 9606 8313 9640 8347
rect 10425 8313 10459 8347
rect 12633 8313 12667 8347
rect 14289 8313 14323 8347
rect 15577 8313 15611 8347
rect 16681 8313 16715 8347
rect 17049 8313 17083 8347
rect 14105 8245 14139 8279
rect 14933 8245 14967 8279
rect 17969 8245 18003 8279
rect 8953 8041 8987 8075
rect 12633 8041 12667 8075
rect 13001 8041 13035 8075
rect 13369 8041 13403 8075
rect 15577 8041 15611 8075
rect 16129 8041 16163 8075
rect 16957 8041 16991 8075
rect 8861 7973 8895 8007
rect 16773 7973 16807 8007
rect 12449 7905 12483 7939
rect 13185 7905 13219 7939
rect 13461 7905 13495 7939
rect 14565 7905 14599 7939
rect 14749 7905 14783 7939
rect 15761 7905 15795 7939
rect 16313 7905 16347 7939
rect 16405 7905 16439 7939
rect 16589 7905 16623 7939
rect 16681 7905 16715 7939
rect 17049 7905 17083 7939
rect 9137 7837 9171 7871
rect 14657 7837 14691 7871
rect 15945 7837 15979 7871
rect 16773 7769 16807 7803
rect 8493 7701 8527 7735
rect 15761 7497 15795 7531
rect 16865 7497 16899 7531
rect 8677 7429 8711 7463
rect 11621 7429 11655 7463
rect 15025 7429 15059 7463
rect 8217 7361 8251 7395
rect 9689 7361 9723 7395
rect 10517 7361 10551 7395
rect 15577 7361 15611 7395
rect 16957 7361 16991 7395
rect 7941 7293 7975 7327
rect 8401 7293 8435 7327
rect 8677 7293 8711 7327
rect 9781 7293 9815 7327
rect 9873 7293 9907 7327
rect 10701 7293 10735 7327
rect 11529 7293 11563 7327
rect 11713 7293 11747 7327
rect 11805 7293 11839 7327
rect 11989 7293 12023 7327
rect 12449 7293 12483 7327
rect 12725 7293 12759 7327
rect 13093 7293 13127 7327
rect 13185 7293 13219 7327
rect 13369 7293 13403 7327
rect 14013 7293 14047 7327
rect 14105 7293 14139 7327
rect 14197 7293 14231 7327
rect 14381 7293 14415 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 15025 7293 15059 7327
rect 15301 7293 15335 7327
rect 15853 7293 15887 7327
rect 16681 7293 16715 7327
rect 6561 7225 6595 7259
rect 10609 7225 10643 7259
rect 12081 7225 12115 7259
rect 12173 7225 12207 7259
rect 12311 7225 12345 7259
rect 12817 7225 12851 7259
rect 12909 7225 12943 7259
rect 13737 7225 13771 7259
rect 15209 7225 15243 7259
rect 8493 7157 8527 7191
rect 10241 7157 10275 7191
rect 11069 7157 11103 7191
rect 12541 7157 12575 7191
rect 13277 7157 13311 7191
rect 14473 7157 14507 7191
rect 14841 7157 14875 7191
rect 15577 7157 15611 7191
rect 16497 7157 16531 7191
rect 9229 6953 9263 6987
rect 10333 6953 10367 6987
rect 12265 6953 12299 6987
rect 12633 6953 12667 6987
rect 12909 6953 12943 6987
rect 13553 6953 13587 6987
rect 8493 6885 8527 6919
rect 9321 6885 9355 6919
rect 10241 6885 10275 6919
rect 14013 6885 14047 6919
rect 15531 6885 15565 6919
rect 8677 6817 8711 6851
rect 8769 6817 8803 6851
rect 10977 6817 11011 6851
rect 11069 6817 11103 6851
rect 11253 6817 11287 6851
rect 12449 6817 12483 6851
rect 12725 6817 12759 6851
rect 12817 6817 12851 6851
rect 13001 6817 13035 6851
rect 13553 6817 13587 6851
rect 13737 6817 13771 6851
rect 13921 6817 13955 6851
rect 14105 6817 14139 6851
rect 14289 6817 14323 6851
rect 14381 6817 14415 6851
rect 14565 6817 14599 6851
rect 15209 6817 15243 6851
rect 15301 6817 15335 6851
rect 15393 6817 15427 6851
rect 16129 6817 16163 6851
rect 9505 6749 9539 6783
rect 10517 6749 10551 6783
rect 15669 6749 15703 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 8861 6681 8895 6715
rect 14565 6681 14599 6715
rect 16313 6681 16347 6715
rect 8493 6613 8527 6647
rect 9873 6613 9907 6647
rect 11253 6613 11287 6647
rect 15025 6613 15059 6647
rect 10241 6341 10275 6375
rect 10609 6341 10643 6375
rect 9873 6205 9907 6239
rect 9965 6205 9999 6239
rect 10241 6205 10275 6239
rect 10333 6205 10367 6239
rect 10425 6205 10459 6239
rect 9606 6137 9640 6171
rect 10609 6137 10643 6171
rect 8493 6069 8527 6103
rect 10057 6069 10091 6103
rect 17040 5797 17074 5831
rect 9321 5729 9355 5763
rect 9588 5729 9622 5763
rect 10977 5729 11011 5763
rect 11244 5729 11278 5763
rect 16773 5729 16807 5763
rect 10701 5525 10735 5559
rect 12357 5525 12391 5559
rect 18153 5525 18187 5559
rect 11161 5185 11195 5219
rect 11417 5117 11451 5151
rect 12541 4981 12575 5015
<< metal1 >>
rect 552 19066 19571 19088
rect 552 19014 5112 19066
rect 5164 19014 5176 19066
rect 5228 19014 5240 19066
rect 5292 19014 5304 19066
rect 5356 19014 5368 19066
rect 5420 19014 9827 19066
rect 9879 19014 9891 19066
rect 9943 19014 9955 19066
rect 10007 19014 10019 19066
rect 10071 19014 10083 19066
rect 10135 19014 14542 19066
rect 14594 19014 14606 19066
rect 14658 19014 14670 19066
rect 14722 19014 14734 19066
rect 14786 19014 14798 19066
rect 14850 19014 19257 19066
rect 19309 19014 19321 19066
rect 19373 19014 19385 19066
rect 19437 19014 19449 19066
rect 19501 19014 19513 19066
rect 19565 19014 19571 19066
rect 552 18992 19571 19014
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 8662 18952 8668 18964
rect 4479 18924 8668 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 9122 18844 9128 18896
rect 9180 18884 9186 18896
rect 9180 18856 9720 18884
rect 9180 18844 9186 18856
rect 842 18776 848 18828
rect 900 18816 906 18828
rect 937 18819 995 18825
rect 937 18816 949 18819
rect 900 18788 949 18816
rect 900 18776 906 18788
rect 937 18785 949 18788
rect 983 18785 995 18819
rect 937 18779 995 18785
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 2593 18819 2651 18825
rect 2593 18816 2605 18819
rect 2556 18788 2605 18816
rect 2556 18776 2562 18788
rect 2593 18785 2605 18788
rect 2639 18785 2651 18819
rect 2593 18779 2651 18785
rect 4154 18776 4160 18828
rect 4212 18816 4218 18828
rect 4249 18819 4307 18825
rect 4249 18816 4261 18819
rect 4212 18788 4261 18816
rect 4212 18776 4218 18788
rect 4249 18785 4261 18788
rect 4295 18785 4307 18819
rect 4249 18779 4307 18785
rect 5810 18776 5816 18828
rect 5868 18816 5874 18828
rect 5905 18819 5963 18825
rect 5905 18816 5917 18819
rect 5868 18788 5917 18816
rect 5868 18776 5874 18788
rect 5905 18785 5917 18788
rect 5951 18785 5963 18819
rect 5905 18779 5963 18785
rect 7466 18776 7472 18828
rect 7524 18816 7530 18828
rect 9692 18825 9720 18856
rect 7561 18819 7619 18825
rect 7561 18816 7573 18819
rect 7524 18788 7573 18816
rect 7524 18776 7530 18788
rect 7561 18785 7573 18788
rect 7607 18785 7619 18819
rect 9217 18819 9275 18825
rect 9217 18816 9229 18819
rect 7561 18779 7619 18785
rect 7668 18788 9229 18816
rect 1213 18751 1271 18757
rect 1213 18717 1225 18751
rect 1259 18748 1271 18751
rect 6454 18748 6460 18760
rect 1259 18720 6460 18748
rect 1259 18717 1271 18720
rect 1213 18711 1271 18717
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 2777 18683 2835 18689
rect 2777 18649 2789 18683
rect 2823 18680 2835 18683
rect 7668 18680 7696 18788
rect 9217 18785 9229 18788
rect 9263 18785 9275 18819
rect 9217 18779 9275 18785
rect 9401 18819 9459 18825
rect 9401 18785 9413 18819
rect 9447 18785 9459 18819
rect 9401 18779 9459 18785
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 9232 18748 9260 18779
rect 9416 18748 9444 18779
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 11149 18819 11207 18825
rect 11149 18816 11161 18819
rect 10836 18788 11161 18816
rect 10836 18776 10842 18788
rect 11149 18785 11161 18788
rect 11195 18785 11207 18819
rect 11149 18779 11207 18785
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 12713 18819 12771 18825
rect 12713 18816 12725 18819
rect 12492 18788 12725 18816
rect 12492 18776 12498 18788
rect 12713 18785 12725 18788
rect 12759 18785 12771 18819
rect 12713 18779 12771 18785
rect 14090 18776 14096 18828
rect 14148 18816 14154 18828
rect 14369 18819 14427 18825
rect 14369 18816 14381 18819
rect 14148 18788 14381 18816
rect 14148 18776 14154 18788
rect 14369 18785 14381 18788
rect 14415 18785 14427 18819
rect 14369 18779 14427 18785
rect 15746 18776 15752 18828
rect 15804 18816 15810 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15804 18788 16313 18816
rect 15804 18776 15810 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 17402 18776 17408 18828
rect 17460 18816 17466 18828
rect 17681 18819 17739 18825
rect 17681 18816 17693 18819
rect 17460 18788 17693 18816
rect 17460 18776 17466 18788
rect 17681 18785 17693 18788
rect 17727 18785 17739 18819
rect 17681 18779 17739 18785
rect 9582 18748 9588 18760
rect 9232 18720 9352 18748
rect 9416 18720 9588 18748
rect 2823 18652 7696 18680
rect 7745 18683 7803 18689
rect 2823 18649 2835 18652
rect 2777 18643 2835 18649
rect 7745 18649 7757 18683
rect 7791 18680 7803 18683
rect 9214 18680 9220 18692
rect 7791 18652 9220 18680
rect 7791 18649 7803 18652
rect 7745 18643 7803 18649
rect 9214 18640 9220 18652
rect 9272 18640 9278 18692
rect 9324 18680 9352 18720
rect 9582 18708 9588 18720
rect 9640 18748 9646 18760
rect 9640 18720 12434 18748
rect 9640 18708 9646 18720
rect 9674 18680 9680 18692
rect 9324 18652 9680 18680
rect 9674 18640 9680 18652
rect 9732 18640 9738 18692
rect 12406 18680 12434 18720
rect 14185 18683 14243 18689
rect 14185 18680 14197 18683
rect 12406 18652 14197 18680
rect 14185 18649 14197 18652
rect 14231 18649 14243 18683
rect 14185 18643 14243 18649
rect 6089 18615 6147 18621
rect 6089 18581 6101 18615
rect 6135 18612 6147 18615
rect 7006 18612 7012 18624
rect 6135 18584 7012 18612
rect 6135 18581 6147 18584
rect 6089 18575 6147 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8570 18572 8576 18624
rect 8628 18612 8634 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 8628 18584 9321 18612
rect 8628 18572 8634 18584
rect 9309 18581 9321 18584
rect 9355 18581 9367 18615
rect 9309 18575 9367 18581
rect 9490 18572 9496 18624
rect 9548 18572 9554 18624
rect 10594 18572 10600 18624
rect 10652 18612 10658 18624
rect 10965 18615 11023 18621
rect 10965 18612 10977 18615
rect 10652 18584 10977 18612
rect 10652 18572 10658 18584
rect 10965 18581 10977 18584
rect 11011 18581 11023 18615
rect 10965 18575 11023 18581
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 16114 18572 16120 18624
rect 16172 18572 16178 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 16816 18584 17509 18612
rect 16816 18572 16822 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 552 18522 19412 18544
rect 552 18470 2755 18522
rect 2807 18470 2819 18522
rect 2871 18470 2883 18522
rect 2935 18470 2947 18522
rect 2999 18470 3011 18522
rect 3063 18470 7470 18522
rect 7522 18470 7534 18522
rect 7586 18470 7598 18522
rect 7650 18470 7662 18522
rect 7714 18470 7726 18522
rect 7778 18470 12185 18522
rect 12237 18470 12249 18522
rect 12301 18470 12313 18522
rect 12365 18470 12377 18522
rect 12429 18470 12441 18522
rect 12493 18470 16900 18522
rect 16952 18470 16964 18522
rect 17016 18470 17028 18522
rect 17080 18470 17092 18522
rect 17144 18470 17156 18522
rect 17208 18470 19412 18522
rect 552 18448 19412 18470
rect 8220 18380 9260 18408
rect 8220 18284 8248 18380
rect 9030 18300 9036 18352
rect 9088 18340 9094 18352
rect 9088 18312 9168 18340
rect 9088 18300 9094 18312
rect 6273 18275 6331 18281
rect 6273 18241 6285 18275
rect 6319 18272 6331 18275
rect 7006 18272 7012 18284
rect 6319 18244 7012 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 8202 18232 8208 18284
rect 8260 18232 8266 18284
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8938 18272 8944 18284
rect 8352 18244 8944 18272
rect 8352 18232 8358 18244
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9140 18281 9168 18312
rect 9125 18275 9183 18281
rect 9125 18241 9137 18275
rect 9171 18241 9183 18275
rect 9232 18272 9260 18380
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 11425 18411 11483 18417
rect 11425 18408 11437 18411
rect 9364 18380 11437 18408
rect 9364 18368 9370 18380
rect 11425 18377 11437 18380
rect 11471 18377 11483 18411
rect 11425 18371 11483 18377
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9232 18244 9873 18272
rect 9125 18235 9183 18241
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 3602 18164 3608 18216
rect 3660 18164 3666 18216
rect 3786 18164 3792 18216
rect 3844 18204 3850 18216
rect 5813 18207 5871 18213
rect 5813 18204 5825 18207
rect 3844 18176 5825 18204
rect 3844 18164 3850 18176
rect 5813 18173 5825 18176
rect 5859 18173 5871 18207
rect 5813 18167 5871 18173
rect 6365 18207 6423 18213
rect 6365 18173 6377 18207
rect 6411 18204 6423 18207
rect 8757 18207 8815 18213
rect 8757 18204 8769 18207
rect 6411 18176 8769 18204
rect 6411 18173 6423 18176
rect 6365 18167 6423 18173
rect 8757 18173 8769 18176
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18204 8907 18207
rect 9398 18204 9404 18216
rect 8895 18176 9404 18204
rect 8895 18173 8907 18176
rect 8849 18167 8907 18173
rect 5568 18139 5626 18145
rect 5568 18105 5580 18139
rect 5614 18136 5626 18139
rect 6089 18139 6147 18145
rect 6089 18136 6101 18139
rect 5614 18108 6101 18136
rect 5614 18105 5626 18108
rect 5568 18099 5626 18105
rect 6089 18105 6101 18108
rect 6135 18105 6147 18139
rect 6089 18099 6147 18105
rect 7960 18139 8018 18145
rect 7960 18105 7972 18139
rect 8006 18136 8018 18139
rect 8294 18136 8300 18148
rect 8006 18108 8300 18136
rect 8006 18105 8018 18108
rect 7960 18099 8018 18105
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 3421 18071 3479 18077
rect 3421 18068 3433 18071
rect 3384 18040 3433 18068
rect 3384 18028 3390 18040
rect 3421 18037 3433 18040
rect 3467 18037 3479 18071
rect 3421 18031 3479 18037
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 4982 18068 4988 18080
rect 4479 18040 4988 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 6730 18028 6736 18080
rect 6788 18028 6794 18080
rect 6822 18028 6828 18080
rect 6880 18028 6886 18080
rect 8386 18028 8392 18080
rect 8444 18028 8450 18080
rect 8772 18068 8800 18167
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18173 9551 18207
rect 9493 18167 9551 18173
rect 8938 18096 8944 18148
rect 8996 18136 9002 18148
rect 9033 18139 9091 18145
rect 9033 18136 9045 18139
rect 8996 18108 9045 18136
rect 8996 18096 9002 18108
rect 9033 18105 9045 18108
rect 9079 18105 9091 18139
rect 9033 18099 9091 18105
rect 9122 18068 9128 18080
rect 8772 18040 9128 18068
rect 9122 18028 9128 18040
rect 9180 18068 9186 18080
rect 9508 18068 9536 18167
rect 9582 18164 9588 18216
rect 9640 18164 9646 18216
rect 11333 18207 11391 18213
rect 11333 18204 11345 18207
rect 11256 18176 11345 18204
rect 9769 18139 9827 18145
rect 9769 18105 9781 18139
rect 9815 18136 9827 18139
rect 10106 18139 10164 18145
rect 10106 18136 10118 18139
rect 9815 18108 10118 18136
rect 9815 18105 9827 18108
rect 9769 18099 9827 18105
rect 10106 18105 10118 18108
rect 10152 18105 10164 18139
rect 10106 18099 10164 18105
rect 11256 18077 11284 18176
rect 11333 18173 11345 18176
rect 11379 18173 11391 18207
rect 11333 18167 11391 18173
rect 16758 18164 16764 18216
rect 16816 18164 16822 18216
rect 9180 18040 9536 18068
rect 11241 18071 11299 18077
rect 9180 18028 9186 18040
rect 11241 18037 11253 18071
rect 11287 18037 11299 18071
rect 11241 18031 11299 18037
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14516 18040 14933 18068
rect 14516 18028 14522 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 16666 18028 16672 18080
rect 16724 18028 16730 18080
rect 552 17978 19571 18000
rect 552 17926 5112 17978
rect 5164 17926 5176 17978
rect 5228 17926 5240 17978
rect 5292 17926 5304 17978
rect 5356 17926 5368 17978
rect 5420 17926 9827 17978
rect 9879 17926 9891 17978
rect 9943 17926 9955 17978
rect 10007 17926 10019 17978
rect 10071 17926 10083 17978
rect 10135 17926 14542 17978
rect 14594 17926 14606 17978
rect 14658 17926 14670 17978
rect 14722 17926 14734 17978
rect 14786 17926 14798 17978
rect 14850 17926 19257 17978
rect 19309 17926 19321 17978
rect 19373 17926 19385 17978
rect 19437 17926 19449 17978
rect 19501 17926 19513 17978
rect 19565 17926 19571 17978
rect 552 17904 19571 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2096 17836 2973 17864
rect 2096 17824 2102 17836
rect 2961 17833 2973 17836
rect 3007 17864 3019 17867
rect 4890 17864 4896 17876
rect 3007 17836 4896 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 6181 17867 6239 17873
rect 6181 17833 6193 17867
rect 6227 17864 6239 17867
rect 6730 17864 6736 17876
rect 6227 17836 6736 17864
rect 6227 17833 6239 17836
rect 6181 17827 6239 17833
rect 6730 17824 6736 17836
rect 6788 17824 6794 17876
rect 8386 17824 8392 17876
rect 8444 17864 8450 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 8444 17836 8493 17864
rect 8444 17824 8450 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 8481 17827 8539 17833
rect 9030 17824 9036 17876
rect 9088 17824 9094 17876
rect 15933 17867 15991 17873
rect 15933 17864 15945 17867
rect 12406 17836 15945 17864
rect 3786 17796 3792 17808
rect 1596 17768 3792 17796
rect 842 17620 848 17672
rect 900 17660 906 17672
rect 1596 17669 1624 17768
rect 1848 17731 1906 17737
rect 1848 17697 1860 17731
rect 1894 17728 1906 17731
rect 2314 17728 2320 17740
rect 1894 17700 2320 17728
rect 1894 17697 1906 17700
rect 1848 17691 1906 17697
rect 2314 17688 2320 17700
rect 2372 17688 2378 17740
rect 3068 17737 3096 17768
rect 3786 17756 3792 17768
rect 3844 17756 3850 17808
rect 3326 17737 3332 17740
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17697 3111 17731
rect 3320 17728 3332 17737
rect 3287 17700 3332 17728
rect 3053 17691 3111 17697
rect 3320 17691 3332 17700
rect 3326 17688 3332 17691
rect 3384 17688 3390 17740
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 5077 17731 5135 17737
rect 5077 17728 5089 17731
rect 4764 17700 5089 17728
rect 4764 17688 4770 17700
rect 5077 17697 5089 17700
rect 5123 17697 5135 17731
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 5077 17691 5135 17697
rect 5460 17700 6745 17728
rect 1581 17663 1639 17669
rect 1581 17660 1593 17663
rect 900 17632 1593 17660
rect 900 17620 906 17632
rect 1581 17629 1593 17632
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 4982 17620 4988 17672
rect 5040 17660 5046 17672
rect 5460 17660 5488 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 7929 17731 7987 17737
rect 7929 17728 7941 17731
rect 6880 17700 7941 17728
rect 6880 17688 6886 17700
rect 7929 17697 7941 17700
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 8386 17688 8392 17740
rect 8444 17728 8450 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 8444 17700 9413 17728
rect 8444 17688 8450 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 5040 17632 5488 17660
rect 5040 17620 5046 17632
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 6512 17632 8217 17660
rect 6512 17620 6518 17632
rect 8205 17629 8217 17632
rect 8251 17660 8263 17663
rect 8294 17660 8300 17672
rect 8251 17632 8300 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 8294 17620 8300 17632
rect 8352 17660 8358 17672
rect 9309 17663 9367 17669
rect 9309 17660 9321 17663
rect 8352 17632 9321 17660
rect 8352 17620 8358 17632
rect 9309 17629 9321 17632
rect 9355 17629 9367 17663
rect 9416 17660 9444 17691
rect 9490 17688 9496 17740
rect 9548 17688 9554 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10226 17728 10232 17740
rect 9732 17700 10232 17728
rect 9732 17688 9738 17700
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 10594 17688 10600 17740
rect 10652 17688 10658 17740
rect 11609 17731 11667 17737
rect 11609 17697 11621 17731
rect 11655 17728 11667 17731
rect 11698 17728 11704 17740
rect 11655 17700 11704 17728
rect 11655 17697 11667 17700
rect 11609 17691 11667 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 12406 17728 12434 17836
rect 15933 17833 15945 17836
rect 15979 17833 15991 17867
rect 15933 17827 15991 17833
rect 14458 17756 14464 17808
rect 14516 17756 14522 17808
rect 16666 17796 16672 17808
rect 15686 17768 16672 17796
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 11756 17700 12434 17728
rect 11756 17688 11762 17700
rect 11422 17660 11428 17672
rect 9416 17632 11428 17660
rect 9309 17623 9367 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 13538 17620 13544 17672
rect 13596 17660 13602 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13596 17632 14197 17660
rect 13596 17620 13602 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 16114 17660 16120 17672
rect 14185 17623 14243 17629
rect 14292 17632 16120 17660
rect 7926 17552 7932 17604
rect 7984 17592 7990 17604
rect 14292 17592 14320 17632
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 7984 17564 14320 17592
rect 7984 17552 7990 17564
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 3292 17496 4445 17524
rect 3292 17484 3298 17496
rect 4433 17493 4445 17496
rect 4479 17524 4491 17527
rect 5258 17524 5264 17536
rect 4479 17496 5264 17524
rect 4479 17493 4491 17496
rect 4433 17487 4491 17493
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5445 17527 5503 17533
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 5626 17524 5632 17536
rect 5491 17496 5632 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 6696 17496 8309 17524
rect 6696 17484 6702 17496
rect 8297 17493 8309 17496
rect 8343 17524 8355 17527
rect 8386 17524 8392 17536
rect 8343 17496 8392 17524
rect 8343 17493 8355 17496
rect 8297 17487 8355 17493
rect 8386 17484 8392 17496
rect 8444 17484 8450 17536
rect 8478 17484 8484 17536
rect 8536 17524 8542 17536
rect 9306 17524 9312 17536
rect 8536 17496 9312 17524
rect 8536 17484 8542 17496
rect 9306 17484 9312 17496
rect 9364 17484 9370 17536
rect 9490 17484 9496 17536
rect 9548 17524 9554 17536
rect 9585 17527 9643 17533
rect 9585 17524 9597 17527
rect 9548 17496 9597 17524
rect 9548 17484 9554 17496
rect 9585 17493 9597 17496
rect 9631 17493 9643 17527
rect 9585 17487 9643 17493
rect 10410 17484 10416 17536
rect 10468 17524 10474 17536
rect 10505 17527 10563 17533
rect 10505 17524 10517 17527
rect 10468 17496 10517 17524
rect 10468 17484 10474 17496
rect 10505 17493 10517 17496
rect 10551 17493 10563 17527
rect 10505 17487 10563 17493
rect 11422 17484 11428 17536
rect 11480 17484 11486 17536
rect 552 17434 19412 17456
rect 552 17382 2755 17434
rect 2807 17382 2819 17434
rect 2871 17382 2883 17434
rect 2935 17382 2947 17434
rect 2999 17382 3011 17434
rect 3063 17382 7470 17434
rect 7522 17382 7534 17434
rect 7586 17382 7598 17434
rect 7650 17382 7662 17434
rect 7714 17382 7726 17434
rect 7778 17382 12185 17434
rect 12237 17382 12249 17434
rect 12301 17382 12313 17434
rect 12365 17382 12377 17434
rect 12429 17382 12441 17434
rect 12493 17382 16900 17434
rect 16952 17382 16964 17434
rect 17016 17382 17028 17434
rect 17080 17382 17092 17434
rect 17144 17382 17156 17434
rect 17208 17382 19412 17434
rect 552 17360 19412 17382
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17320 2467 17323
rect 2685 17323 2743 17329
rect 2685 17320 2697 17323
rect 2455 17292 2697 17320
rect 2455 17289 2467 17292
rect 2409 17283 2467 17289
rect 2685 17289 2697 17292
rect 2731 17289 2743 17323
rect 2685 17283 2743 17289
rect 3513 17323 3571 17329
rect 3513 17289 3525 17323
rect 3559 17320 3571 17323
rect 3602 17320 3608 17332
rect 3559 17292 3608 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 5074 17320 5080 17332
rect 3896 17292 5080 17320
rect 3896 17193 3924 17292
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5534 17280 5540 17332
rect 5592 17320 5598 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 5592 17292 6561 17320
rect 5592 17280 5598 17292
rect 6549 17289 6561 17292
rect 6595 17320 6607 17323
rect 6730 17320 6736 17332
rect 6595 17292 6736 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 6730 17280 6736 17292
rect 6788 17280 6794 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 10781 17323 10839 17329
rect 10781 17320 10793 17323
rect 8904 17292 10793 17320
rect 8904 17280 8910 17292
rect 10781 17289 10793 17292
rect 10827 17289 10839 17323
rect 10781 17283 10839 17289
rect 6822 17252 6828 17264
rect 4448 17224 6828 17252
rect 3881 17187 3939 17193
rect 1780 17156 2176 17184
rect 1780 17125 1808 17156
rect 2148 17128 2176 17156
rect 3881 17153 3893 17187
rect 3927 17184 3939 17187
rect 3970 17184 3976 17196
rect 3927 17156 3976 17184
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 4448 17193 4476 17224
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17184 4767 17187
rect 4755 17156 4936 17184
rect 4755 17153 4767 17156
rect 4709 17147 4767 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1949 17119 2007 17125
rect 1949 17085 1961 17119
rect 1995 17116 2007 17119
rect 2038 17116 2044 17128
rect 1995 17088 2044 17116
rect 1995 17085 2007 17088
rect 1949 17079 2007 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 2130 17076 2136 17128
rect 2188 17116 2194 17128
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 2188 17088 2237 17116
rect 2188 17076 2194 17088
rect 2225 17085 2237 17088
rect 2271 17116 2283 17119
rect 3234 17116 3240 17128
rect 2271 17088 3240 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 3697 17119 3755 17125
rect 3697 17116 3709 17119
rect 3344 17088 3709 17116
rect 3344 17060 3372 17088
rect 3697 17085 3709 17088
rect 3743 17085 3755 17119
rect 3697 17079 3755 17085
rect 4154 17076 4160 17128
rect 4212 17116 4218 17128
rect 4908 17125 4936 17156
rect 5074 17144 5080 17196
rect 5132 17184 5138 17196
rect 5132 17156 6040 17184
rect 5132 17144 5138 17156
rect 4341 17119 4399 17125
rect 4341 17116 4353 17119
rect 4212 17088 4353 17116
rect 4212 17076 4218 17088
rect 4341 17085 4353 17088
rect 4387 17085 4399 17119
rect 4341 17079 4399 17085
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17085 4951 17119
rect 4893 17079 4951 17085
rect 4982 17076 4988 17128
rect 5040 17116 5046 17128
rect 5040 17088 5085 17116
rect 5040 17076 5046 17088
rect 5258 17076 5264 17128
rect 5316 17076 5322 17128
rect 5399 17119 5457 17125
rect 5399 17085 5411 17119
rect 5445 17116 5457 17119
rect 5534 17116 5540 17128
rect 5445 17088 5540 17116
rect 5445 17085 5457 17088
rect 5399 17079 5457 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 5810 17125 5816 17128
rect 5777 17119 5816 17125
rect 5777 17085 5789 17119
rect 5777 17079 5816 17085
rect 5810 17076 5816 17079
rect 5868 17076 5874 17128
rect 6012 17125 6040 17156
rect 5997 17119 6055 17125
rect 5997 17085 6009 17119
rect 6043 17085 6055 17119
rect 5997 17079 6055 17085
rect 6113 17119 6171 17125
rect 6113 17085 6125 17119
rect 6159 17116 6171 17119
rect 6641 17119 6699 17125
rect 6159 17085 6176 17116
rect 6113 17079 6176 17085
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 6687 17088 6776 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 2653 17051 2711 17057
rect 2653 17048 2665 17051
rect 2332 17020 2665 17048
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 2332 16980 2360 17020
rect 2653 17017 2665 17020
rect 2699 17017 2711 17051
rect 2653 17011 2711 17017
rect 2869 17051 2927 17057
rect 2869 17017 2881 17051
rect 2915 17048 2927 17051
rect 3326 17048 3332 17060
rect 2915 17020 3332 17048
rect 2915 17017 2927 17020
rect 2869 17011 2927 17017
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 5169 17051 5227 17057
rect 5169 17017 5181 17051
rect 5215 17017 5227 17051
rect 5169 17011 5227 17017
rect 1903 16952 2360 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 2498 16940 2504 16992
rect 2556 16940 2562 16992
rect 5184 16980 5212 17011
rect 5902 17008 5908 17060
rect 5960 17008 5966 17060
rect 6148 17048 6176 17079
rect 6748 17048 6776 17088
rect 7208 17088 8125 17116
rect 7208 17060 7236 17088
rect 8113 17085 8125 17088
rect 8159 17116 8171 17119
rect 8202 17116 8208 17128
rect 8159 17088 8208 17116
rect 8159 17085 8171 17088
rect 8113 17079 8171 17085
rect 8202 17076 8208 17088
rect 8260 17116 8266 17128
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8260 17088 9229 17116
rect 8260 17076 8266 17088
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 9217 17079 9275 17085
rect 10612 17088 10701 17116
rect 6148 17020 6776 17048
rect 5442 16980 5448 16992
rect 5184 16952 5448 16980
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 5534 16940 5540 16992
rect 5592 16940 5598 16992
rect 5626 16940 5632 16992
rect 5684 16980 5690 16992
rect 6748 16989 6776 17020
rect 7190 17008 7196 17060
rect 7248 17008 7254 17060
rect 7834 17008 7840 17060
rect 7892 17057 7898 17060
rect 7892 17011 7904 17057
rect 9484 17051 9542 17057
rect 9484 17017 9496 17051
rect 9530 17048 9542 17051
rect 9674 17048 9680 17060
rect 9530 17020 9680 17048
rect 9530 17017 9542 17020
rect 9484 17011 9542 17017
rect 7892 17008 7898 17011
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 10612 16989 10640 17088
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 10689 17079 10747 17085
rect 6273 16983 6331 16989
rect 6273 16980 6285 16983
rect 5684 16952 6285 16980
rect 5684 16940 5690 16952
rect 6273 16949 6285 16952
rect 6319 16949 6331 16983
rect 6273 16943 6331 16949
rect 6733 16983 6791 16989
rect 6733 16949 6745 16983
rect 6779 16949 6791 16983
rect 6733 16943 6791 16949
rect 10597 16983 10655 16989
rect 10597 16949 10609 16983
rect 10643 16949 10655 16983
rect 10597 16943 10655 16949
rect 552 16890 19571 16912
rect 552 16838 5112 16890
rect 5164 16838 5176 16890
rect 5228 16838 5240 16890
rect 5292 16838 5304 16890
rect 5356 16838 5368 16890
rect 5420 16838 9827 16890
rect 9879 16838 9891 16890
rect 9943 16838 9955 16890
rect 10007 16838 10019 16890
rect 10071 16838 10083 16890
rect 10135 16838 14542 16890
rect 14594 16838 14606 16890
rect 14658 16838 14670 16890
rect 14722 16838 14734 16890
rect 14786 16838 14798 16890
rect 14850 16838 19257 16890
rect 19309 16838 19321 16890
rect 19373 16838 19385 16890
rect 19437 16838 19449 16890
rect 19501 16838 19513 16890
rect 19565 16838 19571 16890
rect 552 16816 19571 16838
rect 2314 16736 2320 16788
rect 2372 16736 2378 16788
rect 3970 16736 3976 16788
rect 4028 16736 4034 16788
rect 4982 16736 4988 16788
rect 5040 16776 5046 16788
rect 5040 16748 6408 16776
rect 5040 16736 5046 16748
rect 5813 16711 5871 16717
rect 5813 16708 5825 16711
rect 5184 16680 5825 16708
rect 2498 16600 2504 16652
rect 2556 16600 2562 16652
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 5184 16649 5212 16680
rect 5813 16677 5825 16680
rect 5859 16677 5871 16711
rect 6178 16708 6184 16720
rect 5813 16671 5871 16677
rect 6012 16680 6184 16708
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 3292 16612 4077 16640
rect 3292 16600 3298 16612
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 4065 16603 4123 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5534 16640 5540 16652
rect 5399 16612 5540 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5534 16600 5540 16612
rect 5592 16600 5598 16652
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 6012 16649 6040 16680
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 5997 16643 6055 16649
rect 5997 16609 6009 16643
rect 6043 16609 6055 16643
rect 5997 16603 6055 16609
rect 6086 16600 6092 16652
rect 6144 16600 6150 16652
rect 6380 16649 6408 16748
rect 6454 16736 6460 16788
rect 6512 16776 6518 16788
rect 6822 16776 6828 16788
rect 6512 16748 6828 16776
rect 6512 16736 6518 16748
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7101 16779 7159 16785
rect 7101 16745 7113 16779
rect 7147 16776 7159 16779
rect 7193 16779 7251 16785
rect 7193 16776 7205 16779
rect 7147 16748 7205 16776
rect 7147 16745 7159 16748
rect 7101 16739 7159 16745
rect 7193 16745 7205 16748
rect 7239 16745 7251 16779
rect 7193 16739 7251 16745
rect 7834 16736 7840 16788
rect 7892 16736 7898 16788
rect 9033 16779 9091 16785
rect 8220 16748 8984 16776
rect 8220 16708 8248 16748
rect 8754 16708 8760 16720
rect 6932 16680 8248 16708
rect 8312 16680 8760 16708
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 6457 16643 6515 16649
rect 6457 16609 6469 16643
rect 6503 16609 6515 16643
rect 6457 16603 6515 16609
rect 5258 16532 5264 16584
rect 5316 16532 5322 16584
rect 5445 16575 5503 16581
rect 5445 16541 5457 16575
rect 5491 16572 5503 16575
rect 5644 16572 5672 16600
rect 5491 16544 5672 16572
rect 5491 16541 5503 16544
rect 5445 16535 5503 16541
rect 5629 16507 5687 16513
rect 5629 16473 5641 16507
rect 5675 16504 5687 16507
rect 6472 16504 6500 16603
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6696 16612 6745 16640
rect 6696 16600 6702 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 6733 16603 6791 16609
rect 6822 16600 6828 16652
rect 6880 16600 6886 16652
rect 6932 16572 6960 16680
rect 8312 16652 8340 16680
rect 8754 16668 8760 16680
rect 8812 16708 8818 16720
rect 8956 16708 8984 16748
rect 9033 16745 9045 16779
rect 9079 16776 9091 16779
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 9079 16748 9137 16776
rect 9079 16745 9091 16748
rect 9033 16739 9091 16745
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 9732 16748 9781 16776
rect 9732 16736 9738 16748
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 9769 16739 9827 16745
rect 9876 16748 11192 16776
rect 9876 16708 9904 16748
rect 8812 16680 8892 16708
rect 8956 16680 9904 16708
rect 8812 16668 8818 16680
rect 7926 16640 7932 16652
rect 7668 16612 7932 16640
rect 7668 16581 7696 16612
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8294 16600 8300 16652
rect 8352 16600 8358 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 8864 16649 8892 16680
rect 9950 16668 9956 16720
rect 10008 16668 10014 16720
rect 11164 16652 11192 16748
rect 11514 16736 11520 16788
rect 11572 16776 11578 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11572 16748 12081 16776
rect 11572 16736 11578 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 12069 16739 12127 16745
rect 11422 16668 11428 16720
rect 11480 16708 11486 16720
rect 11480 16680 12020 16708
rect 11480 16668 11486 16680
rect 8665 16643 8723 16649
rect 8665 16640 8677 16643
rect 8444 16612 8677 16640
rect 8444 16600 8450 16612
rect 8665 16609 8677 16612
rect 8711 16609 8723 16643
rect 8665 16603 8723 16609
rect 8849 16643 8907 16649
rect 8849 16609 8861 16643
rect 8895 16609 8907 16643
rect 8849 16603 8907 16609
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 9585 16643 9643 16649
rect 9585 16640 9597 16643
rect 9272 16612 9597 16640
rect 9272 16600 9278 16612
rect 9585 16609 9597 16612
rect 9631 16640 9643 16643
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9631 16612 9873 16640
rect 9631 16609 9643 16612
rect 9585 16603 9643 16609
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9861 16603 9919 16609
rect 9968 16612 10057 16640
rect 6656 16544 6960 16572
rect 7561 16575 7619 16581
rect 6656 16513 6684 16544
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 7653 16575 7711 16581
rect 7653 16541 7665 16575
rect 7699 16541 7711 16575
rect 7653 16535 7711 16541
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 5675 16476 6500 16504
rect 6641 16507 6699 16513
rect 5675 16473 5687 16476
rect 5629 16467 5687 16473
rect 6641 16473 6653 16507
rect 6687 16473 6699 16507
rect 6641 16467 6699 16473
rect 7098 16464 7104 16516
rect 7156 16504 7162 16516
rect 7576 16504 7604 16535
rect 8481 16507 8539 16513
rect 8481 16504 8493 16507
rect 7156 16476 8493 16504
rect 7156 16464 7162 16476
rect 8481 16473 8493 16476
rect 8527 16504 8539 16507
rect 9122 16504 9128 16516
rect 8527 16476 9128 16504
rect 8527 16473 8539 16476
rect 8481 16467 8539 16473
rect 9122 16464 9128 16476
rect 9180 16504 9186 16516
rect 9508 16504 9536 16535
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 9968 16572 9996 16612
rect 10045 16609 10057 16612
rect 10091 16640 10103 16643
rect 10226 16640 10232 16652
rect 10091 16612 10232 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 11146 16600 11152 16652
rect 11204 16600 11210 16652
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11790 16640 11796 16652
rect 11296 16612 11796 16640
rect 11296 16600 11302 16612
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 11885 16644 11943 16649
rect 11992 16644 12020 16680
rect 11885 16643 12020 16644
rect 11885 16609 11897 16643
rect 11931 16616 12020 16643
rect 11931 16609 11943 16616
rect 11885 16603 11943 16609
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 12437 16643 12495 16649
rect 12437 16640 12449 16643
rect 12124 16612 12449 16640
rect 12124 16600 12130 16612
rect 12437 16609 12449 16612
rect 12483 16609 12495 16643
rect 12437 16603 12495 16609
rect 9732 16544 9996 16572
rect 11609 16575 11667 16581
rect 9732 16532 9738 16544
rect 11609 16541 11621 16575
rect 11655 16541 11667 16575
rect 11609 16535 11667 16541
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16572 11759 16575
rect 11974 16572 11980 16584
rect 11747 16544 11980 16572
rect 11747 16541 11759 16544
rect 11701 16535 11759 16541
rect 9582 16504 9588 16516
rect 9180 16476 9588 16504
rect 9180 16464 9186 16476
rect 9582 16464 9588 16476
rect 9640 16464 9646 16516
rect 11333 16507 11391 16513
rect 11333 16473 11345 16507
rect 11379 16504 11391 16507
rect 11624 16504 11652 16535
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 12618 16572 12624 16584
rect 12575 16544 12624 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 12268 16504 12296 16535
rect 11379 16476 12296 16504
rect 11379 16473 11391 16476
rect 11333 16467 11391 16473
rect 11808 16448 11836 16476
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 6270 16436 6276 16448
rect 5500 16408 6276 16436
rect 5500 16396 5506 16408
rect 6270 16396 6276 16408
rect 6328 16396 6334 16448
rect 6730 16396 6736 16448
rect 6788 16396 6794 16448
rect 8846 16396 8852 16448
rect 8904 16396 8910 16448
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 10870 16436 10876 16448
rect 8996 16408 10876 16436
rect 8996 16396 9002 16408
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 11425 16439 11483 16445
rect 11425 16405 11437 16439
rect 11471 16436 11483 16439
rect 11606 16436 11612 16448
rect 11471 16408 11612 16436
rect 11471 16405 11483 16408
rect 11425 16399 11483 16405
rect 11606 16396 11612 16408
rect 11664 16396 11670 16448
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 12360 16436 12388 16535
rect 12618 16532 12624 16544
rect 12676 16572 12682 16584
rect 15194 16572 15200 16584
rect 12676 16544 15200 16572
rect 12676 16532 12682 16544
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 12032 16408 12388 16436
rect 12032 16396 12038 16408
rect 552 16346 19412 16368
rect 552 16294 2755 16346
rect 2807 16294 2819 16346
rect 2871 16294 2883 16346
rect 2935 16294 2947 16346
rect 2999 16294 3011 16346
rect 3063 16294 7470 16346
rect 7522 16294 7534 16346
rect 7586 16294 7598 16346
rect 7650 16294 7662 16346
rect 7714 16294 7726 16346
rect 7778 16294 12185 16346
rect 12237 16294 12249 16346
rect 12301 16294 12313 16346
rect 12365 16294 12377 16346
rect 12429 16294 12441 16346
rect 12493 16294 16900 16346
rect 16952 16294 16964 16346
rect 17016 16294 17028 16346
rect 17080 16294 17092 16346
rect 17144 16294 17156 16346
rect 17208 16294 19412 16346
rect 552 16272 19412 16294
rect 4801 16235 4859 16241
rect 4801 16201 4813 16235
rect 4847 16232 4859 16235
rect 5258 16232 5264 16244
rect 4847 16204 5264 16232
rect 4847 16201 4859 16204
rect 4801 16195 4859 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 8478 16232 8484 16244
rect 6328 16204 8484 16232
rect 6328 16192 6334 16204
rect 8478 16192 8484 16204
rect 8536 16192 8542 16244
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9214 16232 9220 16244
rect 8987 16204 9220 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 10502 16232 10508 16244
rect 9324 16204 10508 16232
rect 2130 16124 2136 16176
rect 2188 16124 2194 16176
rect 9324 16164 9352 16204
rect 10502 16192 10508 16204
rect 10560 16232 10566 16244
rect 10560 16204 10824 16232
rect 10560 16192 10566 16204
rect 4540 16136 9352 16164
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2148 16096 2176 16124
rect 4540 16105 4568 16136
rect 9398 16124 9404 16176
rect 9456 16124 9462 16176
rect 9769 16167 9827 16173
rect 9769 16133 9781 16167
rect 9815 16133 9827 16167
rect 9769 16127 9827 16133
rect 1820 16068 2176 16096
rect 4525 16099 4583 16105
rect 1820 16056 1826 16068
rect 2056 16037 2084 16068
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 7098 16056 7104 16108
rect 7156 16056 7162 16108
rect 8754 16056 8760 16108
rect 8812 16056 8818 16108
rect 9784 16096 9812 16127
rect 10796 16105 10824 16204
rect 10870 16192 10876 16244
rect 10928 16232 10934 16244
rect 12526 16232 12532 16244
rect 10928 16204 12532 16232
rect 10928 16192 10934 16204
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 9416 16068 9812 16096
rect 10781 16099 10839 16105
rect 1857 16031 1915 16037
rect 1857 15997 1869 16031
rect 1903 15997 1915 16031
rect 1857 15991 1915 15997
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 1872 15960 1900 15991
rect 2130 15988 2136 16040
rect 2188 15988 2194 16040
rect 2406 15988 2412 16040
rect 2464 16028 2470 16040
rect 2685 16031 2743 16037
rect 2685 16028 2697 16031
rect 2464 16000 2697 16028
rect 2464 15988 2470 16000
rect 2685 15997 2697 16000
rect 2731 16028 2743 16031
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 2731 16000 4445 16028
rect 2731 15997 2743 16000
rect 2685 15991 2743 15997
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 7009 16031 7067 16037
rect 7009 15997 7021 16031
rect 7055 16028 7067 16031
rect 8018 16028 8024 16040
rect 7055 16000 8024 16028
rect 7055 15997 7067 16000
rect 7009 15991 7067 15997
rect 8018 15988 8024 16000
rect 8076 16028 8082 16040
rect 8938 16028 8944 16040
rect 8076 16000 8944 16028
rect 8076 15988 8082 16000
rect 8938 15988 8944 16000
rect 8996 15988 9002 16040
rect 9030 15988 9036 16040
rect 9088 15988 9094 16040
rect 9416 16037 9444 16068
rect 10781 16065 10793 16099
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9582 15988 9588 16040
rect 9640 15988 9646 16040
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10045 16031 10103 16037
rect 9723 16000 9996 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 2222 15960 2228 15972
rect 1872 15932 2228 15960
rect 2222 15920 2228 15932
rect 2280 15920 2286 15972
rect 2498 15920 2504 15972
rect 2556 15920 2562 15972
rect 9600 15960 9628 15988
rect 9769 15963 9827 15969
rect 9769 15960 9781 15963
rect 9600 15932 9781 15960
rect 9769 15929 9781 15932
rect 9815 15929 9827 15963
rect 9968 15960 9996 16000
rect 10045 15997 10057 16031
rect 10091 16028 10103 16031
rect 10594 16028 10600 16040
rect 10091 16000 10600 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10594 15988 10600 16000
rect 10652 15988 10658 16040
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11238 16028 11244 16040
rect 11195 16000 11244 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11238 15988 11244 16000
rect 11296 15988 11302 16040
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 11606 15988 11612 16040
rect 11664 15988 11670 16040
rect 11885 16031 11943 16037
rect 11885 15997 11897 16031
rect 11931 16028 11943 16031
rect 12526 16028 12532 16040
rect 11931 16000 12532 16028
rect 11931 15997 11943 16000
rect 11885 15991 11943 15997
rect 12526 15988 12532 16000
rect 12584 16028 12590 16040
rect 13556 16028 13584 16056
rect 12584 16000 13584 16028
rect 12584 15988 12590 16000
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 10410 15960 10416 15972
rect 9968 15932 10416 15960
rect 9769 15923 9827 15929
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 1302 15852 1308 15904
rect 1360 15892 1366 15904
rect 1673 15895 1731 15901
rect 1673 15892 1685 15895
rect 1360 15864 1685 15892
rect 1360 15852 1366 15864
rect 1673 15861 1685 15864
rect 1719 15861 1731 15895
rect 1673 15855 1731 15861
rect 2869 15895 2927 15901
rect 2869 15861 2881 15895
rect 2915 15892 2927 15895
rect 3234 15892 3240 15904
rect 2915 15864 3240 15892
rect 2915 15861 2927 15864
rect 2869 15855 2927 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 6822 15852 6828 15904
rect 6880 15852 6886 15904
rect 7469 15895 7527 15901
rect 7469 15861 7481 15895
rect 7515 15892 7527 15895
rect 7834 15892 7840 15904
rect 7515 15864 7840 15892
rect 7515 15861 7527 15864
rect 7469 15855 7527 15861
rect 7834 15852 7840 15864
rect 7892 15852 7898 15904
rect 8478 15852 8484 15904
rect 8536 15852 8542 15904
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10229 15895 10287 15901
rect 10229 15892 10241 15895
rect 9999 15864 10241 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10229 15861 10241 15864
rect 10275 15861 10287 15895
rect 11256 15892 11284 15988
rect 11793 15963 11851 15969
rect 11793 15929 11805 15963
rect 11839 15960 11851 15963
rect 12130 15963 12188 15969
rect 12130 15960 12142 15963
rect 11839 15932 12142 15960
rect 11839 15929 11851 15932
rect 11793 15923 11851 15929
rect 12130 15929 12142 15932
rect 12176 15929 12188 15963
rect 12130 15923 12188 15929
rect 12250 15892 12256 15904
rect 11256 15864 12256 15892
rect 10229 15855 10287 15861
rect 12250 15852 12256 15864
rect 12308 15892 12314 15904
rect 13265 15895 13323 15901
rect 13265 15892 13277 15895
rect 12308 15864 13277 15892
rect 12308 15852 12314 15864
rect 13265 15861 13277 15864
rect 13311 15892 13323 15895
rect 14826 15892 14832 15904
rect 13311 15864 14832 15892
rect 13311 15861 13323 15864
rect 13265 15855 13323 15861
rect 14826 15852 14832 15864
rect 14884 15852 14890 15904
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15194 15892 15200 15904
rect 15151 15864 15200 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 552 15802 19571 15824
rect 552 15750 5112 15802
rect 5164 15750 5176 15802
rect 5228 15750 5240 15802
rect 5292 15750 5304 15802
rect 5356 15750 5368 15802
rect 5420 15750 9827 15802
rect 9879 15750 9891 15802
rect 9943 15750 9955 15802
rect 10007 15750 10019 15802
rect 10071 15750 10083 15802
rect 10135 15750 14542 15802
rect 14594 15750 14606 15802
rect 14658 15750 14670 15802
rect 14722 15750 14734 15802
rect 14786 15750 14798 15802
rect 14850 15750 19257 15802
rect 19309 15750 19321 15802
rect 19373 15750 19385 15802
rect 19437 15750 19449 15802
rect 19501 15750 19513 15802
rect 19565 15750 19571 15802
rect 552 15728 19571 15750
rect 1121 15691 1179 15697
rect 1121 15657 1133 15691
rect 1167 15657 1179 15691
rect 1121 15651 1179 15657
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2130 15688 2136 15700
rect 1995 15660 2136 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 845 15555 903 15561
rect 845 15521 857 15555
rect 891 15552 903 15555
rect 1136 15552 1164 15651
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2406 15648 2412 15700
rect 2464 15648 2470 15700
rect 3326 15688 3332 15700
rect 2746 15660 3332 15688
rect 1305 15623 1363 15629
rect 1305 15589 1317 15623
rect 1351 15589 1363 15623
rect 1305 15583 1363 15589
rect 891 15524 1164 15552
rect 891 15521 903 15524
rect 845 15515 903 15521
rect 1320 15416 1348 15583
rect 1762 15580 1768 15632
rect 1820 15580 1826 15632
rect 2041 15623 2099 15629
rect 2041 15589 2053 15623
rect 2087 15620 2099 15623
rect 2222 15620 2228 15632
rect 2087 15592 2228 15620
rect 2087 15589 2099 15592
rect 2041 15583 2099 15589
rect 2222 15580 2228 15592
rect 2280 15580 2286 15632
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2424 15552 2452 15648
rect 2746 15552 2774 15660
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 10502 15648 10508 15700
rect 10560 15648 10566 15700
rect 11330 15648 11336 15700
rect 11388 15648 11394 15700
rect 13081 15691 13139 15697
rect 13081 15657 13093 15691
rect 13127 15688 13139 15691
rect 13814 15688 13820 15700
rect 13127 15660 13820 15688
rect 13127 15657 13139 15660
rect 13081 15651 13139 15657
rect 13814 15648 13820 15660
rect 13872 15648 13878 15700
rect 9398 15629 9404 15632
rect 9392 15620 9404 15629
rect 9359 15592 9404 15620
rect 9392 15583 9404 15592
rect 9398 15580 9404 15583
rect 9456 15580 9462 15632
rect 2179 15524 2452 15552
rect 2608 15524 2774 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 1946 15484 1952 15496
rect 1719 15456 1952 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 1946 15444 1952 15456
rect 2004 15484 2010 15496
rect 2498 15484 2504 15496
rect 2004 15456 2504 15484
rect 2004 15444 2010 15456
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2608 15428 2636 15524
rect 3510 15512 3516 15564
rect 3568 15561 3574 15564
rect 3568 15515 3580 15561
rect 3568 15512 3574 15515
rect 3786 15512 3792 15564
rect 3844 15552 3850 15564
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 3844 15524 6929 15552
rect 3844 15512 3850 15524
rect 6917 15521 6929 15524
rect 6963 15552 6975 15555
rect 7190 15552 7196 15564
rect 6963 15524 7196 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7190 15512 7196 15524
rect 7248 15512 7254 15564
rect 8662 15512 8668 15564
rect 8720 15512 8726 15564
rect 9214 15512 9220 15564
rect 9272 15552 9278 15564
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 9272 15524 10793 15552
rect 9272 15512 9278 15524
rect 10781 15521 10793 15524
rect 10827 15552 10839 15555
rect 10827 15524 11100 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 7208 15484 7236 15512
rect 9122 15484 9128 15496
rect 7208 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 11072 15484 11100 15524
rect 11146 15512 11152 15564
rect 11204 15512 11210 15564
rect 11348 15552 11376 15648
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11348 15524 11437 15552
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 11609 15555 11667 15561
rect 11609 15521 11621 15555
rect 11655 15552 11667 15555
rect 11698 15552 11704 15564
rect 11655 15524 11704 15552
rect 11655 15521 11667 15524
rect 11609 15515 11667 15521
rect 11624 15484 11652 15515
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 11790 15512 11796 15564
rect 11848 15512 11854 15564
rect 11974 15512 11980 15564
rect 12032 15512 12038 15564
rect 12250 15512 12256 15564
rect 12308 15512 12314 15564
rect 12618 15512 12624 15564
rect 12676 15512 12682 15564
rect 12894 15512 12900 15564
rect 12952 15512 12958 15564
rect 11072 15456 11652 15484
rect 10965 15447 11023 15453
rect 2590 15416 2596 15428
rect 1320 15388 2596 15416
rect 2590 15376 2596 15388
rect 2648 15376 2654 15428
rect 10980 15416 11008 15447
rect 11146 15416 11152 15428
rect 10980 15388 11152 15416
rect 11146 15376 11152 15388
rect 11204 15416 11210 15428
rect 11992 15416 12020 15512
rect 11204 15388 12020 15416
rect 11204 15376 11210 15388
rect 1026 15308 1032 15360
rect 1084 15308 1090 15360
rect 1302 15308 1308 15360
rect 1360 15308 1366 15360
rect 2314 15308 2320 15360
rect 2372 15308 2378 15360
rect 10594 15308 10600 15360
rect 10652 15348 10658 15360
rect 10689 15351 10747 15357
rect 10689 15348 10701 15351
rect 10652 15320 10701 15348
rect 10652 15308 10658 15320
rect 10689 15317 10701 15320
rect 10735 15317 10747 15351
rect 10689 15311 10747 15317
rect 11422 15308 11428 15360
rect 11480 15308 11486 15360
rect 11882 15308 11888 15360
rect 11940 15308 11946 15360
rect 552 15258 19412 15280
rect 552 15206 2755 15258
rect 2807 15206 2819 15258
rect 2871 15206 2883 15258
rect 2935 15206 2947 15258
rect 2999 15206 3011 15258
rect 3063 15206 7470 15258
rect 7522 15206 7534 15258
rect 7586 15206 7598 15258
rect 7650 15206 7662 15258
rect 7714 15206 7726 15258
rect 7778 15206 12185 15258
rect 12237 15206 12249 15258
rect 12301 15206 12313 15258
rect 12365 15206 12377 15258
rect 12429 15206 12441 15258
rect 12493 15206 16900 15258
rect 16952 15206 16964 15258
rect 17016 15206 17028 15258
rect 17080 15206 17092 15258
rect 17144 15206 17156 15258
rect 17208 15206 19412 15258
rect 552 15184 19412 15206
rect 2869 15147 2927 15153
rect 2869 15113 2881 15147
rect 2915 15144 2927 15147
rect 3234 15144 3240 15156
rect 2915 15116 3240 15144
rect 2915 15113 2927 15116
rect 2869 15107 2927 15113
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3421 15147 3479 15153
rect 3421 15113 3433 15147
rect 3467 15144 3479 15147
rect 3510 15144 3516 15156
rect 3467 15116 3516 15144
rect 3467 15113 3479 15116
rect 3421 15107 3479 15113
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 8389 15147 8447 15153
rect 8389 15113 8401 15147
rect 8435 15144 8447 15147
rect 9030 15144 9036 15156
rect 8435 15116 9036 15144
rect 8435 15113 8447 15116
rect 8389 15107 8447 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 11514 15104 11520 15156
rect 11572 15104 11578 15156
rect 11701 15147 11759 15153
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 12894 15144 12900 15156
rect 11747 15116 12900 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 3053 15079 3111 15085
rect 3053 15045 3065 15079
rect 3099 15045 3111 15079
rect 3053 15039 3111 15045
rect 842 14968 848 15020
rect 900 14968 906 15020
rect 1112 14943 1170 14949
rect 1112 14909 1124 14943
rect 1158 14909 1170 14943
rect 1112 14903 1170 14909
rect 1026 14832 1032 14884
rect 1084 14872 1090 14884
rect 1136 14872 1164 14903
rect 2314 14900 2320 14952
rect 2372 14940 2378 14952
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 2372 14912 2513 14940
rect 2372 14900 2378 14912
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 3068 14940 3096 15039
rect 3237 14943 3295 14949
rect 3237 14940 3249 14943
rect 3068 14912 3249 14940
rect 2501 14903 2559 14909
rect 3237 14909 3249 14912
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 3605 14943 3663 14949
rect 3605 14909 3617 14943
rect 3651 14909 3663 14943
rect 3605 14903 3663 14909
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 4065 14943 4123 14949
rect 4065 14940 4077 14943
rect 3835 14912 4077 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4065 14909 4077 14912
rect 4111 14940 4123 14943
rect 4154 14940 4160 14952
rect 4111 14912 4160 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 1084 14844 1164 14872
rect 2516 14872 2544 14903
rect 3620 14872 3648 14903
rect 4154 14900 4160 14912
rect 4212 14900 4218 14952
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14940 4307 14943
rect 4798 14940 4804 14952
rect 4295 14912 4804 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 4264 14872 4292 14903
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 4893 14943 4951 14949
rect 4893 14909 4905 14943
rect 4939 14940 4951 14943
rect 5810 14940 5816 14952
rect 4939 14912 5816 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 5810 14900 5816 14912
rect 5868 14900 5874 14952
rect 6270 14900 6276 14952
rect 6328 14900 6334 14952
rect 6540 14943 6598 14949
rect 6540 14909 6552 14943
rect 6586 14940 6598 14943
rect 6822 14940 6828 14952
rect 6586 14912 6828 14940
rect 6586 14909 6598 14912
rect 6540 14903 6598 14909
rect 6822 14900 6828 14912
rect 6880 14900 6886 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9180 14912 9781 14940
rect 9180 14900 9186 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 2516 14844 4292 14872
rect 4433 14875 4491 14881
rect 1084 14832 1090 14844
rect 4433 14841 4445 14875
rect 4479 14872 4491 14875
rect 4522 14872 4528 14884
rect 4479 14844 4528 14872
rect 4479 14841 4491 14844
rect 4433 14835 4491 14841
rect 4522 14832 4528 14844
rect 4580 14872 4586 14884
rect 4709 14875 4767 14881
rect 4709 14872 4721 14875
rect 4580 14844 4721 14872
rect 4580 14832 4586 14844
rect 4709 14841 4721 14844
rect 4755 14841 4767 14875
rect 4709 14835 4767 14841
rect 8938 14832 8944 14884
rect 8996 14872 9002 14884
rect 9502 14875 9560 14881
rect 9502 14872 9514 14875
rect 8996 14844 9514 14872
rect 8996 14832 9002 14844
rect 9502 14841 9514 14844
rect 9548 14841 9560 14875
rect 9502 14835 9560 14841
rect 10594 14832 10600 14884
rect 10652 14872 10658 14884
rect 11606 14881 11612 14884
rect 11333 14875 11391 14881
rect 11333 14872 11345 14875
rect 10652 14844 11345 14872
rect 10652 14832 10658 14844
rect 11333 14841 11345 14844
rect 11379 14841 11391 14875
rect 11333 14835 11391 14841
rect 11549 14875 11612 14881
rect 11549 14841 11561 14875
rect 11595 14841 11612 14875
rect 11549 14835 11612 14841
rect 11606 14832 11612 14835
rect 11664 14872 11670 14884
rect 11882 14872 11888 14884
rect 11664 14844 11888 14872
rect 11664 14832 11670 14844
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 14844 14872 14872 14903
rect 14918 14900 14924 14952
rect 14976 14900 14982 14952
rect 15194 14872 15200 14884
rect 14844 14844 15200 14872
rect 15194 14832 15200 14844
rect 15252 14872 15258 14884
rect 16206 14872 16212 14884
rect 15252 14844 16212 14872
rect 15252 14832 15258 14844
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 2222 14764 2228 14816
rect 2280 14764 2286 14816
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 3973 14807 4031 14813
rect 3973 14773 3985 14807
rect 4019 14804 4031 14807
rect 4154 14804 4160 14816
rect 4019 14776 4160 14804
rect 4019 14773 4031 14776
rect 3973 14767 4031 14773
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 4982 14764 4988 14816
rect 5040 14804 5046 14816
rect 5077 14807 5135 14813
rect 5077 14804 5089 14807
rect 5040 14776 5089 14804
rect 5040 14764 5046 14776
rect 5077 14773 5089 14776
rect 5123 14773 5135 14807
rect 5077 14767 5135 14773
rect 7282 14764 7288 14816
rect 7340 14804 7346 14816
rect 7653 14807 7711 14813
rect 7653 14804 7665 14807
rect 7340 14776 7665 14804
rect 7340 14764 7346 14776
rect 7653 14773 7665 14776
rect 7699 14773 7711 14807
rect 7653 14767 7711 14773
rect 15470 14764 15476 14816
rect 15528 14764 15534 14816
rect 552 14714 19571 14736
rect 552 14662 5112 14714
rect 5164 14662 5176 14714
rect 5228 14662 5240 14714
rect 5292 14662 5304 14714
rect 5356 14662 5368 14714
rect 5420 14662 9827 14714
rect 9879 14662 9891 14714
rect 9943 14662 9955 14714
rect 10007 14662 10019 14714
rect 10071 14662 10083 14714
rect 10135 14662 14542 14714
rect 14594 14662 14606 14714
rect 14658 14662 14670 14714
rect 14722 14662 14734 14714
rect 14786 14662 14798 14714
rect 14850 14662 19257 14714
rect 19309 14662 19321 14714
rect 19373 14662 19385 14714
rect 19437 14662 19449 14714
rect 19501 14662 19513 14714
rect 19565 14662 19571 14714
rect 552 14640 19571 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 3973 14603 4031 14609
rect 1820 14572 2360 14600
rect 1820 14560 1826 14572
rect 2117 14535 2175 14541
rect 2117 14501 2129 14535
rect 2163 14532 2175 14535
rect 2222 14532 2228 14544
rect 2163 14504 2228 14532
rect 2163 14501 2175 14504
rect 2117 14495 2175 14501
rect 2222 14492 2228 14504
rect 2280 14492 2286 14544
rect 2332 14541 2360 14572
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4019 14572 4844 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14501 2375 14535
rect 2317 14495 2375 14501
rect 2866 14492 2872 14544
rect 2924 14532 2930 14544
rect 4062 14532 4068 14544
rect 2924 14504 4068 14532
rect 2924 14492 2930 14504
rect 4062 14492 4068 14504
rect 4120 14532 4126 14544
rect 4157 14535 4215 14541
rect 4157 14532 4169 14535
rect 4120 14504 4169 14532
rect 4120 14492 4126 14504
rect 4157 14501 4169 14504
rect 4203 14501 4215 14535
rect 4157 14495 4215 14501
rect 2240 14396 2268 14492
rect 4522 14424 4528 14476
rect 4580 14424 4586 14476
rect 4816 14473 4844 14572
rect 5810 14560 5816 14612
rect 5868 14560 5874 14612
rect 7834 14560 7840 14612
rect 7892 14560 7898 14612
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14600 8355 14603
rect 8478 14600 8484 14612
rect 8343 14572 8484 14600
rect 8343 14569 8355 14572
rect 8297 14563 8355 14569
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 5074 14492 5080 14544
rect 5132 14532 5138 14544
rect 5261 14535 5319 14541
rect 5261 14532 5273 14535
rect 5132 14504 5273 14532
rect 5132 14492 5138 14504
rect 5261 14501 5273 14504
rect 5307 14532 5319 14535
rect 11422 14532 11428 14544
rect 5307 14504 11428 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 11422 14492 11428 14504
rect 11480 14492 11486 14544
rect 12066 14532 12072 14544
rect 11624 14504 12072 14532
rect 11624 14476 11652 14504
rect 12066 14492 12072 14504
rect 12124 14532 12130 14544
rect 12124 14504 12296 14532
rect 12124 14492 12130 14504
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14433 4859 14467
rect 4801 14427 4859 14433
rect 5534 14424 5540 14476
rect 5592 14464 5598 14476
rect 6926 14467 6984 14473
rect 6926 14464 6938 14467
rect 5592 14436 6938 14464
rect 5592 14424 5598 14436
rect 6926 14433 6938 14436
rect 6972 14433 6984 14467
rect 6926 14427 6984 14433
rect 7098 14424 7104 14476
rect 7156 14424 7162 14476
rect 7190 14424 7196 14476
rect 7248 14424 7254 14476
rect 7282 14424 7288 14476
rect 7340 14424 7346 14476
rect 8757 14467 8815 14473
rect 8757 14464 8769 14467
rect 7576 14436 8769 14464
rect 5442 14396 5448 14408
rect 2240 14368 5448 14396
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 7116 14396 7144 14424
rect 7576 14405 7604 14436
rect 8757 14433 8769 14436
rect 8803 14433 8815 14467
rect 8757 14427 8815 14433
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 11974 14424 11980 14476
rect 12032 14424 12038 14476
rect 12268 14473 12296 14504
rect 15286 14492 15292 14544
rect 15344 14492 15350 14544
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 12084 14436 12173 14464
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7116 14368 7573 14396
rect 7561 14365 7573 14368
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 1946 14288 1952 14340
rect 2004 14288 2010 14340
rect 4893 14331 4951 14337
rect 4893 14297 4905 14331
rect 4939 14328 4951 14331
rect 5166 14328 5172 14340
rect 4939 14300 5172 14328
rect 4939 14297 4951 14300
rect 4893 14291 4951 14297
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 8680 14328 8708 14359
rect 11882 14356 11888 14408
rect 11940 14356 11946 14408
rect 8754 14328 8760 14340
rect 8680 14300 8760 14328
rect 8754 14288 8760 14300
rect 8812 14328 8818 14340
rect 10778 14328 10784 14340
rect 8812 14300 10784 14328
rect 8812 14288 8818 14300
rect 10778 14288 10784 14300
rect 10836 14288 10842 14340
rect 11698 14288 11704 14340
rect 11756 14328 11762 14340
rect 12084 14328 12112 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 12161 14427 12219 14433
rect 12253 14467 12311 14473
rect 12253 14433 12265 14467
rect 12299 14433 12311 14467
rect 12253 14427 12311 14433
rect 12437 14467 12495 14473
rect 12437 14433 12449 14467
rect 12483 14464 12495 14467
rect 12526 14464 12532 14476
rect 12483 14436 12532 14464
rect 12483 14433 12495 14436
rect 12437 14427 12495 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12710 14473 12716 14476
rect 12704 14427 12716 14473
rect 12710 14424 12716 14427
rect 12768 14424 12774 14476
rect 14918 14424 14924 14476
rect 14976 14424 14982 14476
rect 15102 14424 15108 14476
rect 15160 14464 15166 14476
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 15160 14436 15209 14464
rect 15160 14424 15166 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 11756 14300 12112 14328
rect 11756 14288 11762 14300
rect 2130 14220 2136 14272
rect 2188 14220 2194 14272
rect 4154 14220 4160 14272
rect 4212 14220 4218 14272
rect 4614 14220 4620 14272
rect 4672 14220 4678 14272
rect 4982 14220 4988 14272
rect 5040 14260 5046 14272
rect 5261 14263 5319 14269
rect 5261 14260 5273 14263
rect 5040 14232 5273 14260
rect 5040 14220 5046 14232
rect 5261 14229 5273 14232
rect 5307 14229 5319 14263
rect 5261 14223 5319 14229
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 5408 14232 5457 14260
rect 5408 14220 5414 14232
rect 5445 14229 5457 14232
rect 5491 14229 5503 14263
rect 5445 14223 5503 14229
rect 7653 14263 7711 14269
rect 7653 14229 7665 14263
rect 7699 14260 7711 14263
rect 8386 14260 8392 14272
rect 7699 14232 8392 14260
rect 7699 14229 7711 14232
rect 7653 14223 7711 14229
rect 8386 14220 8392 14232
rect 8444 14220 8450 14272
rect 11606 14220 11612 14272
rect 11664 14220 11670 14272
rect 11977 14263 12035 14269
rect 11977 14229 11989 14263
rect 12023 14260 12035 14263
rect 12802 14260 12808 14272
rect 12023 14232 12808 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13814 14220 13820 14272
rect 13872 14220 13878 14272
rect 552 14170 19412 14192
rect 552 14118 2755 14170
rect 2807 14118 2819 14170
rect 2871 14118 2883 14170
rect 2935 14118 2947 14170
rect 2999 14118 3011 14170
rect 3063 14118 7470 14170
rect 7522 14118 7534 14170
rect 7586 14118 7598 14170
rect 7650 14118 7662 14170
rect 7714 14118 7726 14170
rect 7778 14118 12185 14170
rect 12237 14118 12249 14170
rect 12301 14118 12313 14170
rect 12365 14118 12377 14170
rect 12429 14118 12441 14170
rect 12493 14118 16900 14170
rect 16952 14118 16964 14170
rect 17016 14118 17028 14170
rect 17080 14118 17092 14170
rect 17144 14118 17156 14170
rect 17208 14118 19412 14170
rect 552 14096 19412 14118
rect 3329 14059 3387 14065
rect 3329 14025 3341 14059
rect 3375 14056 3387 14059
rect 4338 14056 4344 14068
rect 3375 14028 4344 14056
rect 3375 14025 3387 14028
rect 3329 14019 3387 14025
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4985 14059 5043 14065
rect 4724 14028 4936 14056
rect 2774 13920 2780 13932
rect 1872 13892 2780 13920
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 1872 13861 1900 13892
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 4724 13929 4752 14028
rect 4798 13948 4804 14000
rect 4856 13948 4862 14000
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 4709 13883 4767 13889
rect 1673 13855 1731 13861
rect 1673 13852 1685 13855
rect 1360 13824 1685 13852
rect 1360 13812 1366 13824
rect 1673 13821 1685 13824
rect 1719 13821 1731 13855
rect 1673 13815 1731 13821
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2179 13824 2360 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2332 13728 2360 13824
rect 2958 13812 2964 13864
rect 3016 13812 3022 13864
rect 4453 13855 4511 13861
rect 4453 13821 4465 13855
rect 4499 13852 4511 13855
rect 4614 13852 4620 13864
rect 4499 13824 4620 13852
rect 4499 13821 4511 13824
rect 4453 13815 4511 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4816 13852 4844 13948
rect 4908 13920 4936 14028
rect 4985 14025 4997 14059
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5000 13988 5028 14019
rect 5534 14016 5540 14068
rect 5592 14016 5598 14068
rect 11241 14059 11299 14065
rect 11241 14025 11253 14059
rect 11287 14056 11299 14059
rect 11698 14056 11704 14068
rect 11287 14028 11704 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12529 14059 12587 14065
rect 12529 14056 12541 14059
rect 12124 14028 12541 14056
rect 12124 14016 12130 14028
rect 12529 14025 12541 14028
rect 12575 14025 12587 14059
rect 12529 14019 12587 14025
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12768 14028 12909 14056
rect 12768 14016 12774 14028
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 5810 13988 5816 14000
rect 5000 13960 5816 13988
rect 5810 13948 5816 13960
rect 5868 13948 5874 14000
rect 7282 13988 7288 14000
rect 6656 13960 7288 13988
rect 5626 13920 5632 13932
rect 4908 13892 5632 13920
rect 5626 13880 5632 13892
rect 5684 13920 5690 13932
rect 6270 13920 6276 13932
rect 5684 13892 6276 13920
rect 5684 13880 5690 13892
rect 6270 13880 6276 13892
rect 6328 13880 6334 13932
rect 6656 13929 6684 13960
rect 7282 13948 7288 13960
rect 7340 13948 7346 14000
rect 11425 13991 11483 13997
rect 11425 13988 11437 13991
rect 10980 13960 11437 13988
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6914 13880 6920 13932
rect 6972 13880 6978 13932
rect 4816 13824 5028 13852
rect 4338 13744 4344 13796
rect 4396 13784 4402 13796
rect 4801 13787 4859 13793
rect 4801 13784 4813 13787
rect 4396 13756 4813 13784
rect 4396 13744 4402 13756
rect 4801 13753 4813 13756
rect 4847 13753 4859 13787
rect 4801 13747 4859 13753
rect 2314 13676 2320 13728
rect 2372 13676 2378 13728
rect 5000 13725 5028 13824
rect 5350 13812 5356 13864
rect 5408 13812 5414 13864
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 5500 13824 6561 13852
rect 5500 13812 5506 13824
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 8444 13824 9873 13852
rect 8444 13812 8450 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10091 13824 10885 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10873 13821 10885 13824
rect 10919 13852 10931 13855
rect 10980 13852 11008 13960
rect 11425 13957 11437 13960
rect 11471 13957 11483 13991
rect 11716 13988 11744 14016
rect 13909 13991 13967 13997
rect 13909 13988 13921 13991
rect 11716 13960 12388 13988
rect 11425 13951 11483 13957
rect 10919 13824 11008 13852
rect 11149 13855 11207 13861
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11882 13852 11888 13864
rect 11195 13824 11888 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11882 13812 11888 13824
rect 11940 13852 11946 13864
rect 12176 13861 12204 13960
rect 12360 13920 12388 13960
rect 12452 13960 13921 13988
rect 12452 13929 12480 13960
rect 13909 13957 13921 13960
rect 13955 13957 13967 13991
rect 13909 13951 13967 13957
rect 12437 13923 12495 13929
rect 12437 13920 12449 13923
rect 12360 13892 12449 13920
rect 12437 13889 12449 13892
rect 12483 13889 12495 13923
rect 12437 13883 12495 13889
rect 12161 13855 12219 13861
rect 11940 13824 12112 13852
rect 11940 13812 11946 13824
rect 11054 13744 11060 13796
rect 11112 13744 11118 13796
rect 11425 13787 11483 13793
rect 11425 13753 11437 13787
rect 11471 13784 11483 13787
rect 11514 13784 11520 13796
rect 11471 13756 11520 13784
rect 11471 13753 11483 13756
rect 11425 13747 11483 13753
rect 11514 13744 11520 13756
rect 11572 13744 11578 13796
rect 12084 13784 12112 13824
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12618 13852 12624 13864
rect 12161 13815 12219 13821
rect 12268 13824 12624 13852
rect 12268 13784 12296 13824
rect 12618 13812 12624 13824
rect 12676 13812 12682 13864
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 12802 13852 12808 13864
rect 12759 13824 12808 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13872 13824 14013 13852
rect 13872 13812 13878 13824
rect 14001 13821 14013 13824
rect 14047 13852 14059 13855
rect 15102 13852 15108 13864
rect 14047 13824 15108 13852
rect 14047 13821 14059 13824
rect 14001 13815 14059 13821
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 16206 13812 16212 13864
rect 16264 13812 16270 13864
rect 16482 13812 16488 13864
rect 16540 13812 16546 13864
rect 12084 13756 12296 13784
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 5000 13719 5059 13725
rect 5000 13688 5013 13719
rect 5001 13685 5013 13688
rect 5047 13685 5059 13719
rect 5001 13679 5059 13685
rect 5166 13676 5172 13728
rect 5224 13716 5230 13728
rect 5442 13716 5448 13728
rect 5224 13688 5448 13716
rect 5224 13676 5230 13688
rect 5442 13676 5448 13688
rect 5500 13676 5506 13728
rect 9953 13719 10011 13725
rect 9953 13685 9965 13719
rect 9999 13716 10011 13719
rect 10226 13716 10232 13728
rect 9999 13688 10232 13716
rect 9999 13685 10011 13688
rect 9953 13679 10011 13685
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 10689 13719 10747 13725
rect 10689 13685 10701 13719
rect 10735 13716 10747 13719
rect 10870 13716 10876 13728
rect 10735 13688 10876 13716
rect 10735 13685 10747 13688
rect 10689 13679 10747 13685
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11701 13719 11759 13725
rect 11701 13685 11713 13719
rect 11747 13716 11759 13719
rect 11790 13716 11796 13728
rect 11747 13688 11796 13716
rect 11747 13685 11759 13688
rect 11701 13679 11759 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 552 13626 19571 13648
rect 552 13574 5112 13626
rect 5164 13574 5176 13626
rect 5228 13574 5240 13626
rect 5292 13574 5304 13626
rect 5356 13574 5368 13626
rect 5420 13574 9827 13626
rect 9879 13574 9891 13626
rect 9943 13574 9955 13626
rect 10007 13574 10019 13626
rect 10071 13574 10083 13626
rect 10135 13574 14542 13626
rect 14594 13574 14606 13626
rect 14658 13574 14670 13626
rect 14722 13574 14734 13626
rect 14786 13574 14798 13626
rect 14850 13574 19257 13626
rect 19309 13574 19321 13626
rect 19373 13574 19385 13626
rect 19437 13574 19449 13626
rect 19501 13574 19513 13626
rect 19565 13574 19571 13626
rect 552 13552 19571 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2593 13515 2651 13521
rect 2593 13512 2605 13515
rect 2372 13484 2605 13512
rect 2372 13472 2378 13484
rect 2593 13481 2605 13484
rect 2639 13481 2651 13515
rect 2593 13475 2651 13481
rect 5074 13472 5080 13524
rect 5132 13472 5138 13524
rect 7745 13515 7803 13521
rect 7745 13481 7757 13515
rect 7791 13512 7803 13515
rect 11146 13512 11152 13524
rect 7791 13484 11152 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 11701 13515 11759 13521
rect 11701 13481 11713 13515
rect 11747 13481 11759 13515
rect 15010 13512 15016 13524
rect 11701 13475 11759 13481
rect 14936 13484 15016 13512
rect 1302 13453 1308 13456
rect 1296 13444 1308 13453
rect 1263 13416 1308 13444
rect 1296 13407 1308 13416
rect 1302 13404 1308 13407
rect 1360 13404 1366 13456
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 4985 13447 5043 13453
rect 4985 13444 4997 13447
rect 4120 13416 4997 13444
rect 4120 13404 4126 13416
rect 4985 13413 4997 13416
rect 5031 13413 5043 13447
rect 5092 13444 5120 13472
rect 5169 13447 5227 13453
rect 5169 13444 5181 13447
rect 5092 13416 5181 13444
rect 4985 13407 5043 13413
rect 5169 13413 5181 13416
rect 5215 13413 5227 13447
rect 5169 13407 5227 13413
rect 7834 13404 7840 13456
rect 7892 13444 7898 13456
rect 8573 13447 8631 13453
rect 8573 13444 8585 13447
rect 7892 13416 8585 13444
rect 7892 13404 7898 13416
rect 8573 13413 8585 13416
rect 8619 13413 8631 13447
rect 8573 13407 8631 13413
rect 8757 13447 8815 13453
rect 8757 13413 8769 13447
rect 8803 13444 8815 13447
rect 9030 13444 9036 13456
rect 8803 13416 9036 13444
rect 8803 13413 8815 13416
rect 8757 13407 8815 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 11716 13444 11744 13475
rect 12314 13447 12372 13453
rect 12314 13444 12326 13447
rect 9456 13416 11652 13444
rect 11716 13416 12326 13444
rect 9456 13404 9462 13416
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 2498 13376 2504 13388
rect 2096 13348 2504 13376
rect 2096 13336 2102 13348
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 2774 13336 2780 13388
rect 2832 13336 2838 13388
rect 2961 13379 3019 13385
rect 2961 13345 2973 13379
rect 3007 13376 3019 13379
rect 3142 13376 3148 13388
rect 3007 13348 3148 13376
rect 3007 13345 3019 13348
rect 2961 13339 3019 13345
rect 3142 13336 3148 13348
rect 3200 13376 3206 13388
rect 4080 13376 4108 13404
rect 3200 13348 4108 13376
rect 3200 13336 3206 13348
rect 5442 13336 5448 13388
rect 5500 13376 5506 13388
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 5500 13348 6009 13376
rect 5500 13336 5506 13348
rect 5997 13345 6009 13348
rect 6043 13345 6055 13379
rect 5997 13339 6055 13345
rect 6914 13336 6920 13388
rect 6972 13376 6978 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 6972 13348 7481 13376
rect 6972 13336 6978 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 8389 13379 8447 13385
rect 8389 13376 8401 13379
rect 8067 13348 8401 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 8389 13345 8401 13348
rect 8435 13345 8447 13379
rect 8389 13339 8447 13345
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 9309 13379 9367 13385
rect 9309 13376 9321 13379
rect 9180 13348 9321 13376
rect 9180 13336 9186 13348
rect 9309 13345 9321 13348
rect 9355 13345 9367 13379
rect 9309 13339 9367 13345
rect 9576 13379 9634 13385
rect 9576 13345 9588 13379
rect 9622 13376 9634 13379
rect 9950 13376 9956 13388
rect 9622 13348 9956 13376
rect 9622 13345 9634 13348
rect 9576 13339 9634 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 1029 13311 1087 13317
rect 1029 13277 1041 13311
rect 1075 13277 1087 13311
rect 1029 13271 1087 13277
rect 1044 13172 1072 13271
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 4764 13280 5825 13308
rect 4764 13268 4770 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 5813 13271 5871 13277
rect 5920 13280 7665 13308
rect 4430 13200 4436 13252
rect 4488 13240 4494 13252
rect 5920 13240 5948 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 8294 13268 8300 13320
rect 8352 13268 8358 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13277 11575 13311
rect 11624 13308 11652 13416
rect 12314 13413 12326 13416
rect 12360 13413 12372 13447
rect 12314 13407 12372 13413
rect 11698 13336 11704 13388
rect 11756 13336 11762 13388
rect 11790 13336 11796 13388
rect 11848 13336 11854 13388
rect 11974 13336 11980 13388
rect 12032 13336 12038 13388
rect 14936 13385 14964 13484
rect 15010 13472 15016 13484
rect 15068 13512 15074 13524
rect 16482 13512 16488 13524
rect 15068 13484 16488 13512
rect 15068 13472 15074 13484
rect 16482 13472 16488 13484
rect 16540 13472 16546 13524
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13345 14979 13379
rect 14921 13339 14979 13345
rect 15102 13336 15108 13388
rect 15160 13336 15166 13388
rect 16206 13336 16212 13388
rect 16264 13336 16270 13388
rect 16482 13336 16488 13388
rect 16540 13376 16546 13388
rect 16577 13379 16635 13385
rect 16577 13376 16589 13379
rect 16540 13348 16589 13376
rect 16540 13336 16546 13348
rect 16577 13345 16589 13348
rect 16623 13345 16635 13379
rect 16577 13339 16635 13345
rect 11992 13308 12020 13336
rect 11624 13280 12020 13308
rect 11517 13271 11575 13277
rect 4488 13212 5948 13240
rect 10689 13243 10747 13249
rect 4488 13200 4494 13212
rect 10689 13209 10701 13243
rect 10735 13240 10747 13243
rect 11330 13240 11336 13252
rect 10735 13212 11336 13240
rect 10735 13209 10747 13212
rect 10689 13203 10747 13209
rect 11330 13200 11336 13212
rect 11388 13240 11394 13252
rect 11532 13240 11560 13271
rect 12066 13268 12072 13320
rect 12124 13268 12130 13320
rect 15289 13243 15347 13249
rect 15289 13240 15301 13243
rect 11388 13212 11560 13240
rect 15212 13212 15301 13240
rect 11388 13200 11394 13212
rect 15212 13184 15240 13212
rect 15289 13209 15301 13212
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 1762 13172 1768 13184
rect 1044 13144 1768 13172
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 2958 13172 2964 13184
rect 2455 13144 2964 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 2958 13132 2964 13144
rect 3016 13172 3022 13184
rect 3970 13172 3976 13184
rect 3016 13144 3976 13172
rect 3016 13132 3022 13144
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 6086 13132 6092 13184
rect 6144 13172 6150 13184
rect 6181 13175 6239 13181
rect 6181 13172 6193 13175
rect 6144 13144 6193 13172
rect 6144 13132 6150 13144
rect 6181 13141 6193 13144
rect 6227 13141 6239 13175
rect 6181 13135 6239 13141
rect 10962 13132 10968 13184
rect 11020 13132 11026 13184
rect 13449 13175 13507 13181
rect 13449 13141 13461 13175
rect 13495 13172 13507 13175
rect 13722 13172 13728 13184
rect 13495 13144 13728 13172
rect 13495 13141 13507 13144
rect 13449 13135 13507 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 15194 13132 15200 13184
rect 15252 13132 15258 13184
rect 17862 13132 17868 13184
rect 17920 13132 17926 13184
rect 552 13082 19412 13104
rect 552 13030 2755 13082
rect 2807 13030 2819 13082
rect 2871 13030 2883 13082
rect 2935 13030 2947 13082
rect 2999 13030 3011 13082
rect 3063 13030 7470 13082
rect 7522 13030 7534 13082
rect 7586 13030 7598 13082
rect 7650 13030 7662 13082
rect 7714 13030 7726 13082
rect 7778 13030 12185 13082
rect 12237 13030 12249 13082
rect 12301 13030 12313 13082
rect 12365 13030 12377 13082
rect 12429 13030 12441 13082
rect 12493 13030 16900 13082
rect 16952 13030 16964 13082
rect 17016 13030 17028 13082
rect 17080 13030 17092 13082
rect 17144 13030 17156 13082
rect 17208 13030 19412 13082
rect 552 13008 19412 13030
rect 2774 12928 2780 12980
rect 2832 12968 2838 12980
rect 3973 12971 4031 12977
rect 3973 12968 3985 12971
rect 2832 12940 3985 12968
rect 2832 12928 2838 12940
rect 3973 12937 3985 12940
rect 4019 12937 4031 12971
rect 3973 12931 4031 12937
rect 4430 12928 4436 12980
rect 4488 12928 4494 12980
rect 5626 12928 5632 12980
rect 5684 12928 5690 12980
rect 8021 12971 8079 12977
rect 8021 12937 8033 12971
rect 8067 12968 8079 12971
rect 8294 12968 8300 12980
rect 8067 12940 8300 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 9674 12968 9680 12980
rect 8588 12940 9680 12968
rect 8110 12860 8116 12912
rect 8168 12900 8174 12912
rect 8588 12900 8616 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9950 12928 9956 12980
rect 10008 12928 10014 12980
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 10367 12940 11008 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 8168 12872 8616 12900
rect 8168 12860 8174 12872
rect 8662 12860 8668 12912
rect 8720 12900 8726 12912
rect 9493 12903 9551 12909
rect 9493 12900 9505 12903
rect 8720 12872 9505 12900
rect 8720 12860 8726 12872
rect 9493 12869 9505 12872
rect 9539 12869 9551 12903
rect 9493 12863 9551 12869
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 10781 12903 10839 12909
rect 10781 12900 10793 12903
rect 10744 12872 10793 12900
rect 10744 12860 10750 12872
rect 10781 12869 10793 12872
rect 10827 12869 10839 12903
rect 10980 12900 11008 12940
rect 11054 12928 11060 12980
rect 11112 12968 11118 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 11112 12940 11253 12968
rect 11112 12928 11118 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12526 12968 12532 12980
rect 12124 12940 12532 12968
rect 12124 12928 12130 12940
rect 12526 12928 12532 12940
rect 12584 12968 12590 12980
rect 12805 12971 12863 12977
rect 12805 12968 12817 12971
rect 12584 12940 12817 12968
rect 12584 12928 12590 12940
rect 12805 12937 12817 12940
rect 12851 12937 12863 12971
rect 12805 12931 12863 12937
rect 11698 12900 11704 12912
rect 10980 12872 11704 12900
rect 10781 12863 10839 12869
rect 11698 12860 11704 12872
rect 11756 12860 11762 12912
rect 2498 12792 2504 12844
rect 2556 12832 2562 12844
rect 2556 12804 2728 12832
rect 2556 12792 2562 12804
rect 1213 12767 1271 12773
rect 1213 12733 1225 12767
rect 1259 12764 1271 12767
rect 1762 12764 1768 12776
rect 1259 12736 1768 12764
rect 1259 12733 1271 12736
rect 1213 12727 1271 12733
rect 1762 12724 1768 12736
rect 1820 12764 1826 12776
rect 2590 12764 2596 12776
rect 1820 12736 2596 12764
rect 1820 12724 1826 12736
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 2700 12773 2728 12804
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 9030 12832 9036 12844
rect 8128 12804 9036 12832
rect 2685 12767 2743 12773
rect 2685 12733 2697 12767
rect 2731 12733 2743 12767
rect 2685 12727 2743 12733
rect 2866 12724 2872 12776
rect 2924 12724 2930 12776
rect 3789 12767 3847 12773
rect 3789 12764 3801 12767
rect 3068 12736 3801 12764
rect 1480 12699 1538 12705
rect 1480 12665 1492 12699
rect 1526 12696 1538 12699
rect 2777 12699 2835 12705
rect 2777 12696 2789 12699
rect 1526 12668 2789 12696
rect 1526 12665 1538 12668
rect 1480 12659 1538 12665
rect 2777 12665 2789 12668
rect 2823 12665 2835 12699
rect 2777 12659 2835 12665
rect 2593 12631 2651 12637
rect 2593 12597 2605 12631
rect 2639 12628 2651 12631
rect 2682 12628 2688 12640
rect 2639 12600 2688 12628
rect 2639 12597 2651 12600
rect 2593 12591 2651 12597
rect 2682 12588 2688 12600
rect 2740 12628 2746 12640
rect 3068 12628 3096 12736
rect 3789 12733 3801 12736
rect 3835 12764 3847 12767
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 3835 12736 4169 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12733 4307 12767
rect 4724 12764 4752 12792
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4724 12736 4905 12764
rect 4249 12727 4307 12733
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 3970 12656 3976 12708
rect 4028 12656 4034 12708
rect 2740 12600 3096 12628
rect 2740 12588 2746 12600
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 3237 12631 3295 12637
rect 3237 12628 3249 12631
rect 3200 12600 3249 12628
rect 3200 12588 3206 12600
rect 3237 12597 3249 12600
rect 3283 12597 3295 12631
rect 4264 12628 4292 12727
rect 5442 12724 5448 12776
rect 5500 12724 5506 12776
rect 6914 12724 6920 12776
rect 6972 12724 6978 12776
rect 7190 12724 7196 12776
rect 7248 12724 7254 12776
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8128 12773 8156 12804
rect 9030 12792 9036 12804
rect 9088 12792 9094 12844
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10962 12832 10968 12844
rect 10459 12804 10968 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10962 12792 10968 12804
rect 11020 12792 11026 12844
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7892 12736 7941 12764
rect 7892 12724 7898 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8113 12767 8171 12773
rect 8113 12733 8125 12767
rect 8159 12733 8171 12767
rect 8113 12727 8171 12733
rect 8386 12724 8392 12776
rect 8444 12724 8450 12776
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9398 12764 9404 12776
rect 8996 12736 9404 12764
rect 8996 12724 9002 12736
rect 9398 12724 9404 12736
rect 9456 12764 9462 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9456 12736 9505 12764
rect 9456 12724 9462 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 9769 12767 9827 12773
rect 9769 12764 9781 12767
rect 9732 12736 9781 12764
rect 9732 12724 9738 12736
rect 9769 12733 9781 12736
rect 9815 12733 9827 12767
rect 9769 12727 9827 12733
rect 10137 12767 10195 12773
rect 10137 12733 10149 12767
rect 10183 12764 10195 12767
rect 10226 12764 10232 12776
rect 10183 12736 10232 12764
rect 10183 12733 10195 12736
rect 10137 12727 10195 12733
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10318 12724 10324 12776
rect 10376 12764 10382 12776
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 10376 12736 10517 12764
rect 10376 12724 10382 12736
rect 10505 12733 10517 12736
rect 10551 12764 10563 12767
rect 10551 12736 10732 12764
rect 10551 12733 10563 12736
rect 10505 12727 10563 12733
rect 4614 12656 4620 12708
rect 4672 12696 4678 12708
rect 4709 12699 4767 12705
rect 4709 12696 4721 12699
rect 4672 12668 4721 12696
rect 4672 12656 4678 12668
rect 4709 12665 4721 12668
rect 4755 12696 4767 12699
rect 5460 12696 5488 12724
rect 4755 12668 5488 12696
rect 8404 12696 8432 12724
rect 8404 12668 9444 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 9416 12640 9444 12668
rect 4890 12628 4896 12640
rect 4264 12600 4896 12628
rect 3237 12591 3295 12597
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5442 12628 5448 12640
rect 5123 12600 5448 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7098 12628 7104 12640
rect 7055 12600 7104 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 8938 12628 8944 12640
rect 8619 12600 8944 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 9398 12588 9404 12640
rect 9456 12588 9462 12640
rect 9677 12631 9735 12637
rect 9677 12597 9689 12631
rect 9723 12628 9735 12631
rect 10226 12628 10232 12640
rect 9723 12600 10232 12628
rect 9723 12597 9735 12600
rect 9677 12591 9735 12597
rect 10226 12588 10232 12600
rect 10284 12628 10290 12640
rect 10597 12631 10655 12637
rect 10597 12628 10609 12631
rect 10284 12600 10609 12628
rect 10284 12588 10290 12600
rect 10597 12597 10609 12600
rect 10643 12597 10655 12631
rect 10704 12628 10732 12736
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10928 12736 11069 12764
rect 10928 12724 10934 12736
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 11330 12724 11336 12776
rect 11388 12724 11394 12776
rect 14185 12767 14243 12773
rect 14185 12733 14197 12767
rect 14231 12764 14243 12767
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14231 12736 14841 12764
rect 14231 12733 14243 12736
rect 14185 12727 14243 12733
rect 14829 12733 14841 12736
rect 14875 12764 14887 12767
rect 15010 12764 15016 12776
rect 14875 12736 15016 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15102 12724 15108 12776
rect 15160 12724 15166 12776
rect 10781 12699 10839 12705
rect 10781 12665 10793 12699
rect 10827 12696 10839 12699
rect 10962 12696 10968 12708
rect 10827 12668 10968 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 11020 12668 11468 12696
rect 11020 12656 11026 12668
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10704 12600 10885 12628
rect 10597 12591 10655 12597
rect 10873 12597 10885 12600
rect 10919 12597 10931 12631
rect 11440 12628 11468 12668
rect 11514 12656 11520 12708
rect 11572 12656 11578 12708
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 13633 12699 13691 12705
rect 13633 12696 13645 12699
rect 13412 12668 13645 12696
rect 13412 12656 13418 12668
rect 13633 12665 13645 12668
rect 13679 12665 13691 12699
rect 16298 12696 16304 12708
rect 15962 12668 16304 12696
rect 13633 12659 13691 12665
rect 16298 12656 16304 12668
rect 16356 12656 16362 12708
rect 13372 12628 13400 12656
rect 11440 12600 13400 12628
rect 10873 12591 10931 12597
rect 552 12538 19571 12560
rect 552 12486 5112 12538
rect 5164 12486 5176 12538
rect 5228 12486 5240 12538
rect 5292 12486 5304 12538
rect 5356 12486 5368 12538
rect 5420 12486 9827 12538
rect 9879 12486 9891 12538
rect 9943 12486 9955 12538
rect 10007 12486 10019 12538
rect 10071 12486 10083 12538
rect 10135 12486 14542 12538
rect 14594 12486 14606 12538
rect 14658 12486 14670 12538
rect 14722 12486 14734 12538
rect 14786 12486 14798 12538
rect 14850 12486 19257 12538
rect 19309 12486 19321 12538
rect 19373 12486 19385 12538
rect 19437 12486 19449 12538
rect 19501 12486 19513 12538
rect 19565 12486 19571 12538
rect 552 12464 19571 12486
rect 2406 12384 2412 12436
rect 2464 12384 2470 12436
rect 2572 12427 2630 12433
rect 2572 12424 2584 12427
rect 2516 12396 2584 12424
rect 2516 12300 2544 12396
rect 2572 12393 2584 12396
rect 2618 12393 2630 12427
rect 2572 12387 2630 12393
rect 2866 12384 2872 12436
rect 2924 12384 2930 12436
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5445 12427 5503 12433
rect 5445 12424 5457 12427
rect 5040 12396 5457 12424
rect 5040 12384 5046 12396
rect 5445 12393 5457 12396
rect 5491 12393 5503 12427
rect 5813 12427 5871 12433
rect 5813 12424 5825 12427
rect 5445 12387 5503 12393
rect 5552 12396 5825 12424
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 3234 12356 3240 12368
rect 2832 12328 3240 12356
rect 2832 12316 2838 12328
rect 3234 12316 3240 12328
rect 3292 12316 3298 12368
rect 2498 12248 2504 12300
rect 2556 12248 2562 12300
rect 3142 12248 3148 12300
rect 3200 12248 3206 12300
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4246 12288 4252 12300
rect 4203 12260 4252 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 4246 12248 4252 12260
rect 4304 12248 4310 12300
rect 4614 12248 4620 12300
rect 4672 12248 4678 12300
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 5552 12288 5580 12396
rect 5813 12393 5825 12396
rect 5859 12393 5871 12427
rect 10962 12424 10968 12436
rect 5813 12387 5871 12393
rect 10428 12396 10968 12424
rect 5626 12316 5632 12368
rect 5684 12356 5690 12368
rect 5684 12328 7236 12356
rect 5684 12316 5690 12328
rect 4856 12260 5580 12288
rect 6937 12291 6995 12297
rect 4856 12248 4862 12260
rect 6937 12257 6949 12291
rect 6983 12288 6995 12291
rect 7098 12288 7104 12300
rect 6983 12260 7104 12288
rect 6983 12257 6995 12260
rect 6937 12251 6995 12257
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7208 12297 7236 12328
rect 10134 12316 10140 12368
rect 10192 12356 10198 12368
rect 10428 12356 10456 12396
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12676 12396 12725 12424
rect 12676 12384 12682 12396
rect 12713 12393 12725 12396
rect 12759 12393 12771 12427
rect 12713 12387 12771 12393
rect 12066 12356 12072 12368
rect 10192 12328 10456 12356
rect 10192 12316 10198 12328
rect 7193 12291 7251 12297
rect 7193 12257 7205 12291
rect 7239 12288 7251 12291
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7239 12260 7757 12288
rect 7239 12257 7251 12260
rect 7193 12251 7251 12257
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 7745 12251 7803 12257
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 10428 12297 10456 12328
rect 10980 12328 12072 12356
rect 10980 12297 11008 12328
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 14001 12359 14059 12365
rect 14001 12325 14013 12359
rect 14047 12356 14059 12359
rect 14458 12356 14464 12368
rect 14047 12328 14464 12356
rect 14047 12325 14059 12328
rect 14001 12319 14059 12325
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 14921 12359 14979 12365
rect 14921 12325 14933 12359
rect 14967 12356 14979 12359
rect 15010 12356 15016 12368
rect 14967 12328 15016 12356
rect 14967 12325 14979 12328
rect 14921 12319 14979 12325
rect 15010 12316 15016 12328
rect 15068 12316 15074 12368
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 9456 12260 10333 12288
rect 9456 12248 9462 12260
rect 10321 12257 10333 12260
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 10413 12291 10471 12297
rect 10413 12257 10425 12291
rect 10459 12257 10471 12291
rect 10413 12251 10471 12257
rect 10965 12291 11023 12297
rect 10965 12257 10977 12291
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11221 12291 11279 12297
rect 11221 12288 11233 12291
rect 11112 12260 11233 12288
rect 11112 12248 11118 12260
rect 11221 12257 11233 12260
rect 11267 12257 11279 12291
rect 11221 12251 11279 12257
rect 12805 12291 12863 12297
rect 12805 12257 12817 12291
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12220 2927 12223
rect 3050 12220 3056 12232
rect 2915 12192 3056 12220
rect 2915 12189 2927 12192
rect 2869 12183 2927 12189
rect 3050 12180 3056 12192
rect 3108 12220 3114 12232
rect 3326 12220 3332 12232
rect 3108 12192 3332 12220
rect 3108 12180 3114 12192
rect 3326 12180 3332 12192
rect 3384 12180 3390 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 4890 12180 4896 12232
rect 4948 12180 4954 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 6086 12220 6092 12232
rect 5123 12192 6092 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 8021 12223 8079 12229
rect 8021 12189 8033 12223
rect 8067 12220 8079 12223
rect 8478 12220 8484 12232
rect 8067 12192 8484 12220
rect 8067 12189 8079 12192
rect 8021 12183 8079 12189
rect 8478 12180 8484 12192
rect 8536 12180 8542 12232
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12220 9367 12223
rect 9766 12220 9772 12232
rect 9355 12192 9772 12220
rect 9355 12189 9367 12192
rect 9309 12183 9367 12189
rect 9766 12180 9772 12192
rect 9824 12220 9830 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9824 12192 10057 12220
rect 9824 12180 9830 12192
rect 10045 12189 10057 12192
rect 10091 12220 10103 12223
rect 10226 12220 10232 12232
rect 10091 12192 10232 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 10226 12180 10232 12192
rect 10284 12220 10290 12232
rect 10505 12223 10563 12229
rect 10505 12220 10517 12223
rect 10284 12192 10517 12220
rect 10284 12180 10290 12192
rect 10505 12189 10517 12192
rect 10551 12189 10563 12223
rect 10505 12183 10563 12189
rect 10597 12223 10655 12229
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10870 12220 10876 12232
rect 10643 12192 10876 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 5629 12155 5687 12161
rect 5629 12121 5641 12155
rect 5675 12152 5687 12155
rect 5675 12124 6316 12152
rect 5675 12121 5687 12124
rect 5629 12115 5687 12121
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12084 2651 12087
rect 2682 12084 2688 12096
rect 2639 12056 2688 12084
rect 2639 12053 2651 12056
rect 2593 12047 2651 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3053 12087 3111 12093
rect 3053 12053 3065 12087
rect 3099 12084 3111 12087
rect 3142 12084 3148 12096
rect 3099 12056 3148 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4433 12087 4491 12093
rect 4433 12084 4445 12087
rect 4120 12056 4445 12084
rect 4120 12044 4126 12056
rect 4433 12053 4445 12056
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 5442 12044 5448 12096
rect 5500 12044 5506 12096
rect 6288 12084 6316 12124
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10612 12152 10640 12183
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 12820 12220 12848 12251
rect 13354 12248 13360 12300
rect 13412 12248 13418 12300
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13722 12288 13728 12300
rect 13679 12260 13728 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13648 12220 13676 12251
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14093 12291 14151 12297
rect 14093 12257 14105 12291
rect 14139 12257 14151 12291
rect 14093 12251 14151 12257
rect 12820 12192 13676 12220
rect 9916 12124 10640 12152
rect 12345 12155 12403 12161
rect 9916 12112 9922 12124
rect 12345 12121 12357 12155
rect 12391 12152 12403 12155
rect 14108 12152 14136 12251
rect 12391 12124 14136 12152
rect 12391 12121 12403 12124
rect 12345 12115 12403 12121
rect 7190 12084 7196 12096
rect 6288 12056 7196 12084
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 9490 12044 9496 12096
rect 9548 12044 9554 12096
rect 10781 12087 10839 12093
rect 10781 12053 10793 12087
rect 10827 12084 10839 12087
rect 10870 12084 10876 12096
rect 10827 12056 10876 12084
rect 10827 12053 10839 12056
rect 10781 12047 10839 12053
rect 10870 12044 10876 12056
rect 10928 12044 10934 12096
rect 552 11994 19412 12016
rect 552 11942 2755 11994
rect 2807 11942 2819 11994
rect 2871 11942 2883 11994
rect 2935 11942 2947 11994
rect 2999 11942 3011 11994
rect 3063 11942 7470 11994
rect 7522 11942 7534 11994
rect 7586 11942 7598 11994
rect 7650 11942 7662 11994
rect 7714 11942 7726 11994
rect 7778 11942 12185 11994
rect 12237 11942 12249 11994
rect 12301 11942 12313 11994
rect 12365 11942 12377 11994
rect 12429 11942 12441 11994
rect 12493 11942 16900 11994
rect 16952 11942 16964 11994
rect 17016 11942 17028 11994
rect 17080 11942 17092 11994
rect 17144 11942 17156 11994
rect 17208 11942 19412 11994
rect 552 11920 19412 11942
rect 2685 11883 2743 11889
rect 2685 11849 2697 11883
rect 2731 11880 2743 11883
rect 3142 11880 3148 11892
rect 2731 11852 3148 11880
rect 2731 11849 2743 11852
rect 2685 11843 2743 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 4890 11840 4896 11892
rect 4948 11840 4954 11892
rect 5169 11883 5227 11889
rect 5169 11849 5181 11883
rect 5215 11880 5227 11883
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5215 11852 5457 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 5445 11843 5503 11849
rect 5920 11852 7665 11880
rect 4706 11772 4712 11824
rect 4764 11812 4770 11824
rect 5920 11812 5948 11852
rect 7653 11849 7665 11852
rect 7699 11880 7711 11883
rect 7834 11880 7840 11892
rect 7699 11852 7840 11880
rect 7699 11849 7711 11852
rect 7653 11843 7711 11849
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 10873 11883 10931 11889
rect 10873 11849 10885 11883
rect 10919 11880 10931 11883
rect 11054 11880 11060 11892
rect 10919 11852 11060 11880
rect 10919 11849 10931 11852
rect 10873 11843 10931 11849
rect 11054 11840 11060 11852
rect 11112 11840 11118 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15378 11880 15384 11892
rect 15252 11852 15384 11880
rect 15252 11840 15258 11852
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 15930 11840 15936 11892
rect 15988 11880 15994 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15988 11852 16221 11880
rect 15988 11840 15994 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 16209 11843 16267 11849
rect 4764 11784 5948 11812
rect 4764 11772 4770 11784
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2958 11744 2964 11756
rect 2363 11716 2964 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2958 11704 2964 11716
rect 3016 11744 3022 11756
rect 3234 11744 3240 11756
rect 3016 11716 3240 11744
rect 3016 11704 3022 11716
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 5626 11744 5632 11756
rect 5552 11716 5632 11744
rect 2498 11636 2504 11688
rect 2556 11636 2562 11688
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3513 11679 3571 11685
rect 3513 11676 3525 11679
rect 2648 11648 3525 11676
rect 2648 11636 2654 11648
rect 3513 11645 3525 11648
rect 3559 11676 3571 11679
rect 5552 11676 5580 11716
rect 5626 11704 5632 11716
rect 5684 11744 5690 11756
rect 5810 11744 5816 11756
rect 5684 11716 5816 11744
rect 5684 11704 5690 11716
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5920 11685 5948 11784
rect 13446 11772 13452 11824
rect 13504 11812 13510 11824
rect 16666 11812 16672 11824
rect 13504 11784 16672 11812
rect 13504 11772 13510 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 6273 11747 6331 11753
rect 6273 11713 6285 11747
rect 6319 11713 6331 11747
rect 6273 11707 6331 11713
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 3559 11648 5580 11676
rect 5644 11648 5917 11676
rect 3559 11645 3571 11648
rect 3513 11639 3571 11645
rect 2516 11608 2544 11636
rect 3050 11608 3056 11620
rect 2516 11580 3056 11608
rect 3050 11568 3056 11580
rect 3108 11568 3114 11620
rect 3780 11611 3838 11617
rect 3780 11577 3792 11611
rect 3826 11608 3838 11611
rect 3970 11608 3976 11620
rect 3826 11580 3976 11608
rect 3826 11577 3838 11580
rect 3780 11571 3838 11577
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 5644 11617 5672 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6086 11636 6092 11688
rect 6144 11636 6150 11688
rect 4985 11611 5043 11617
rect 4985 11577 4997 11611
rect 5031 11577 5043 11611
rect 4985 11571 5043 11577
rect 5201 11611 5259 11617
rect 5201 11577 5213 11611
rect 5247 11608 5259 11611
rect 5629 11611 5687 11617
rect 5247 11580 5580 11608
rect 5247 11577 5259 11580
rect 5201 11571 5259 11577
rect 3326 11500 3332 11552
rect 3384 11540 3390 11552
rect 5000 11540 5028 11571
rect 3384 11512 5028 11540
rect 5353 11543 5411 11549
rect 3384 11500 3390 11512
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 5442 11540 5448 11552
rect 5399 11512 5448 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 5552 11540 5580 11580
rect 5629 11577 5641 11611
rect 5675 11577 5687 11611
rect 5629 11571 5687 11577
rect 5813 11611 5871 11617
rect 5813 11577 5825 11611
rect 5859 11608 5871 11611
rect 6104 11608 6132 11636
rect 5859 11580 6132 11608
rect 5859 11577 5871 11580
rect 5813 11571 5871 11577
rect 5905 11543 5963 11549
rect 5905 11540 5917 11543
rect 5552 11512 5917 11540
rect 5905 11509 5917 11512
rect 5951 11509 5963 11543
rect 5905 11503 5963 11509
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6288 11540 6316 11707
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 10134 11744 10140 11756
rect 8444 11716 10140 11744
rect 8444 11704 8450 11716
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 15746 11744 15752 11756
rect 14516 11716 15752 11744
rect 14516 11704 14522 11716
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 16758 11744 16764 11756
rect 15804 11716 16764 11744
rect 15804 11704 15810 11716
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 13728 11688 13780 11694
rect 8294 11636 8300 11688
rect 8352 11676 8358 11688
rect 9766 11676 9772 11688
rect 8352 11648 9772 11676
rect 8352 11636 8358 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 10594 11636 10600 11688
rect 10652 11636 10658 11688
rect 10686 11636 10692 11688
rect 10744 11636 10750 11688
rect 10870 11636 10876 11688
rect 10928 11636 10934 11688
rect 12618 11636 12624 11688
rect 12676 11676 12682 11688
rect 13354 11676 13360 11688
rect 12676 11648 13360 11676
rect 12676 11636 12682 11648
rect 13354 11636 13360 11648
rect 13412 11676 13418 11688
rect 13633 11679 13691 11685
rect 13633 11676 13645 11679
rect 13412 11648 13645 11676
rect 13412 11636 13418 11648
rect 13633 11645 13645 11648
rect 13679 11645 13691 11679
rect 13633 11639 13691 11645
rect 15194 11636 15200 11688
rect 15252 11636 15258 11688
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15381 11679 15439 11685
rect 15381 11676 15393 11679
rect 15344 11648 15393 11676
rect 15344 11636 15350 11648
rect 15381 11645 15393 11648
rect 15427 11676 15439 11679
rect 16022 11676 16028 11688
rect 15427 11648 16028 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 16022 11636 16028 11648
rect 16080 11676 16086 11688
rect 16117 11679 16175 11685
rect 16117 11676 16129 11679
rect 16080 11648 16129 11676
rect 16080 11636 16086 11648
rect 16117 11645 16129 11648
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 16393 11679 16451 11685
rect 16393 11676 16405 11679
rect 16356 11648 16405 11676
rect 16356 11636 16362 11648
rect 16393 11645 16405 11648
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 13728 11630 13780 11636
rect 6540 11611 6598 11617
rect 6540 11577 6552 11611
rect 6586 11608 6598 11611
rect 6638 11608 6644 11620
rect 6586 11580 6644 11608
rect 6586 11577 6598 11580
rect 6540 11571 6598 11577
rect 6638 11568 6644 11580
rect 6696 11568 6702 11620
rect 8846 11568 8852 11620
rect 8904 11608 8910 11620
rect 9858 11608 9864 11620
rect 8904 11580 9864 11608
rect 8904 11568 8910 11580
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 14182 11568 14188 11620
rect 14240 11608 14246 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 14240 11580 14381 11608
rect 14240 11568 14246 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 14369 11571 14427 11577
rect 14918 11568 14924 11620
rect 14976 11608 14982 11620
rect 15304 11608 15332 11636
rect 14976 11580 15332 11608
rect 14976 11568 14982 11580
rect 6052 11512 6316 11540
rect 9309 11543 9367 11549
rect 6052 11500 6058 11512
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9582 11540 9588 11552
rect 9355 11512 9588 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10410 11500 10416 11552
rect 10468 11540 10474 11552
rect 10594 11540 10600 11552
rect 10468 11512 10600 11540
rect 10468 11500 10474 11512
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 15286 11500 15292 11552
rect 15344 11500 15350 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 16390 11540 16396 11552
rect 15528 11512 16396 11540
rect 15528 11500 15534 11512
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 16669 11543 16727 11549
rect 16669 11509 16681 11543
rect 16715 11540 16727 11543
rect 16850 11540 16856 11552
rect 16715 11512 16856 11540
rect 16715 11509 16727 11512
rect 16669 11503 16727 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 552 11450 19571 11472
rect 552 11398 5112 11450
rect 5164 11398 5176 11450
rect 5228 11398 5240 11450
rect 5292 11398 5304 11450
rect 5356 11398 5368 11450
rect 5420 11398 9827 11450
rect 9879 11398 9891 11450
rect 9943 11398 9955 11450
rect 10007 11398 10019 11450
rect 10071 11398 10083 11450
rect 10135 11398 14542 11450
rect 14594 11398 14606 11450
rect 14658 11398 14670 11450
rect 14722 11398 14734 11450
rect 14786 11398 14798 11450
rect 14850 11398 19257 11450
rect 19309 11398 19321 11450
rect 19373 11398 19385 11450
rect 19437 11398 19449 11450
rect 19501 11398 19513 11450
rect 19565 11398 19571 11450
rect 552 11376 19571 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11305 2191 11339
rect 2133 11299 2191 11305
rect 2041 11203 2099 11209
rect 2041 11169 2053 11203
rect 2087 11200 2099 11203
rect 2148 11200 2176 11299
rect 3142 11296 3148 11348
rect 3200 11296 3206 11348
rect 4062 11296 4068 11348
rect 4120 11296 4126 11348
rect 4246 11296 4252 11348
rect 4304 11296 4310 11348
rect 4693 11339 4751 11345
rect 4693 11305 4705 11339
rect 4739 11336 4751 11339
rect 6086 11336 6092 11348
rect 4739 11308 6092 11336
rect 4739 11305 4751 11308
rect 4693 11299 4751 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6638 11296 6644 11348
rect 6696 11296 6702 11348
rect 8205 11339 8263 11345
rect 8205 11305 8217 11339
rect 8251 11336 8263 11339
rect 8386 11336 8392 11348
rect 8251 11308 8392 11336
rect 8251 11305 8263 11308
rect 8205 11299 8263 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 9766 11336 9772 11348
rect 8588 11308 9772 11336
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 2777 11271 2835 11277
rect 2777 11268 2789 11271
rect 2363 11240 2789 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 2777 11237 2789 11240
rect 2823 11237 2835 11271
rect 3160 11268 3188 11296
rect 2777 11231 2835 11237
rect 2884 11240 3188 11268
rect 2087 11172 2176 11200
rect 2685 11203 2743 11209
rect 2087 11169 2099 11172
rect 2041 11163 2099 11169
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 2884 11200 2912 11240
rect 4798 11228 4804 11280
rect 4856 11268 4862 11280
rect 4893 11271 4951 11277
rect 4893 11268 4905 11271
rect 4856 11240 4905 11268
rect 4856 11228 4862 11240
rect 4893 11237 4905 11240
rect 4939 11237 4951 11271
rect 4893 11231 4951 11237
rect 8294 11228 8300 11280
rect 8352 11228 8358 11280
rect 2731 11172 2912 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 2958 11160 2964 11212
rect 3016 11160 3022 11212
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3145 11203 3203 11209
rect 3145 11200 3157 11203
rect 3108 11172 3157 11200
rect 3108 11160 3114 11172
rect 3145 11169 3157 11172
rect 3191 11200 3203 11203
rect 3697 11203 3755 11209
rect 3697 11200 3709 11203
rect 3191 11172 3709 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3697 11169 3709 11172
rect 3743 11169 3755 11203
rect 3697 11163 3755 11169
rect 2976 11132 3004 11160
rect 2976 11104 3188 11132
rect 3160 11076 3188 11104
rect 3142 11024 3148 11076
rect 3200 11024 3206 11076
rect 3712 11064 3740 11163
rect 5442 11160 5448 11212
rect 5500 11200 5506 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 5500 11172 6469 11200
rect 5500 11160 5506 11172
rect 6457 11169 6469 11172
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11200 8447 11203
rect 8588 11200 8616 11308
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10226 11345 10232 11348
rect 10045 11339 10103 11345
rect 10045 11305 10057 11339
rect 10091 11305 10103 11339
rect 10045 11299 10103 11305
rect 10203 11339 10232 11345
rect 10203 11305 10215 11339
rect 10203 11299 10232 11305
rect 9490 11268 9496 11280
rect 8956 11240 9496 11268
rect 8435 11172 8616 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8846 11160 8852 11212
rect 8904 11160 8910 11212
rect 8956 11209 8984 11240
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 10060 11268 10088 11299
rect 10226 11296 10232 11299
rect 10284 11296 10290 11348
rect 15841 11339 15899 11345
rect 14016 11308 15700 11336
rect 9600 11240 10088 11268
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9600 11200 9628 11240
rect 10410 11228 10416 11280
rect 10468 11228 10474 11280
rect 13078 11268 13084 11280
rect 12834 11240 13084 11268
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 9263 11172 9628 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9674 11160 9680 11212
rect 9732 11160 9738 11212
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10318 11200 10324 11212
rect 9824 11172 10324 11200
rect 9824 11160 9830 11172
rect 10318 11160 10324 11172
rect 10376 11160 10382 11212
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11885 11203 11943 11209
rect 11885 11200 11897 11203
rect 11388 11172 11897 11200
rect 11388 11160 11394 11172
rect 11885 11169 11897 11172
rect 11931 11169 11943 11203
rect 11885 11163 11943 11169
rect 12618 11160 12624 11212
rect 12676 11160 12682 11212
rect 13354 11160 13360 11212
rect 13412 11200 13418 11212
rect 14016 11209 14044 11308
rect 15286 11268 15292 11280
rect 14660 11240 15292 11268
rect 14001 11203 14059 11209
rect 14001 11200 14013 11203
rect 13412 11172 14013 11200
rect 13412 11160 13418 11172
rect 14001 11169 14013 11172
rect 14047 11169 14059 11203
rect 14001 11163 14059 11169
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 14660 11209 14688 11240
rect 15286 11228 15292 11240
rect 15344 11228 15350 11280
rect 15672 11212 15700 11308
rect 15841 11305 15853 11339
rect 15887 11336 15899 11339
rect 15930 11336 15936 11348
rect 15887 11308 15936 11336
rect 15887 11305 15899 11308
rect 15841 11299 15899 11305
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 16482 11336 16488 11348
rect 16080 11308 16488 11336
rect 16080 11296 16086 11308
rect 16482 11296 16488 11308
rect 16540 11296 16546 11348
rect 15948 11268 15976 11296
rect 15948 11240 16436 11268
rect 14645 11203 14703 11209
rect 14645 11169 14657 11203
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 14734 11160 14740 11212
rect 14792 11160 14798 11212
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11169 14887 11203
rect 14947 11203 15005 11209
rect 14947 11200 14959 11203
rect 14829 11163 14887 11169
rect 14936 11169 14959 11200
rect 14993 11169 15005 11203
rect 14936 11163 15005 11169
rect 8021 11135 8079 11141
rect 8021 11101 8033 11135
rect 8067 11132 8079 11135
rect 9490 11132 9496 11144
rect 8067 11104 9496 11132
rect 8067 11101 8079 11104
rect 8021 11095 8079 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 11422 11132 11428 11144
rect 9631 11104 11428 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14844 11132 14872 11163
rect 14516 11104 14872 11132
rect 14516 11092 14522 11104
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 3712 11036 4537 11064
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 4525 11027 4583 11033
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 9953 11067 10011 11073
rect 8343 11036 9260 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 1854 10956 1860 11008
rect 1912 10956 1918 11008
rect 2317 10999 2375 11005
rect 2317 10965 2329 10999
rect 2363 10996 2375 10999
rect 3326 10996 3332 11008
rect 2363 10968 3332 10996
rect 2363 10965 2375 10968
rect 2317 10959 2375 10965
rect 3326 10956 3332 10968
rect 3384 10996 3390 11008
rect 4065 10999 4123 11005
rect 4065 10996 4077 10999
rect 3384 10968 4077 10996
rect 3384 10956 3390 10968
rect 4065 10965 4077 10968
rect 4111 10965 4123 10999
rect 4065 10959 4123 10965
rect 4709 10999 4767 11005
rect 4709 10965 4721 10999
rect 4755 10996 4767 10999
rect 4890 10996 4896 11008
rect 4755 10968 4896 10996
rect 4755 10965 4767 10968
rect 4709 10959 4767 10965
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 9030 10956 9036 11008
rect 9088 10956 9094 11008
rect 9232 10996 9260 11036
rect 9953 11033 9965 11067
rect 9999 11064 10011 11067
rect 10134 11064 10140 11076
rect 9999 11036 10140 11064
rect 9999 11033 10011 11036
rect 9953 11027 10011 11033
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 14001 11067 14059 11073
rect 14001 11064 14013 11067
rect 13872 11036 14013 11064
rect 13872 11024 13878 11036
rect 14001 11033 14013 11036
rect 14047 11064 14059 11067
rect 14936 11064 14964 11163
rect 15102 11160 15108 11212
rect 15160 11200 15166 11212
rect 15470 11200 15476 11212
rect 15160 11172 15476 11200
rect 15160 11160 15166 11172
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15654 11160 15660 11212
rect 15712 11160 15718 11212
rect 15746 11160 15752 11212
rect 15804 11160 15810 11212
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11200 15991 11203
rect 16022 11200 16028 11212
rect 15979 11172 16028 11200
rect 15979 11169 15991 11172
rect 15933 11163 15991 11169
rect 16022 11160 16028 11172
rect 16080 11160 16086 11212
rect 16298 11160 16304 11212
rect 16356 11160 16362 11212
rect 16408 11209 16436 11240
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11169 16451 11203
rect 16393 11163 16451 11169
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 16577 11163 16635 11169
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 16592 11132 16620 11163
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16724 11172 16773 11200
rect 16724 11160 16730 11172
rect 16761 11169 16773 11172
rect 16807 11169 16819 11203
rect 16761 11163 16819 11169
rect 16850 11160 16856 11212
rect 16908 11160 16914 11212
rect 16945 11203 17003 11209
rect 16945 11169 16957 11203
rect 16991 11169 17003 11203
rect 16945 11163 17003 11169
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17218 11200 17224 11212
rect 17175 11172 17224 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 16960 11132 16988 11163
rect 17218 11160 17224 11172
rect 17276 11160 17282 11212
rect 15611 11104 16988 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 16117 11067 16175 11073
rect 16117 11064 16129 11067
rect 14047 11036 14964 11064
rect 15120 11036 16129 11064
rect 14047 11033 14059 11036
rect 14001 11027 14059 11033
rect 15120 11008 15148 11036
rect 16117 11033 16129 11036
rect 16163 11033 16175 11067
rect 16117 11027 16175 11033
rect 16390 11024 16396 11076
rect 16448 11064 16454 11076
rect 16485 11067 16543 11073
rect 16485 11064 16497 11067
rect 16448 11036 16497 11064
rect 16448 11024 16454 11036
rect 16485 11033 16497 11036
rect 16531 11033 16543 11067
rect 17129 11067 17187 11073
rect 17129 11064 17141 11067
rect 16485 11027 16543 11033
rect 16592 11036 17141 11064
rect 10229 10999 10287 11005
rect 10229 10996 10241 10999
rect 9232 10968 10241 10996
rect 10229 10965 10241 10968
rect 10275 10965 10287 10999
rect 10229 10959 10287 10965
rect 14458 10956 14464 11008
rect 14516 10956 14522 11008
rect 15102 10956 15108 11008
rect 15160 10956 15166 11008
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 15562 10996 15568 11008
rect 15344 10968 15568 10996
rect 15344 10956 15350 10968
rect 15562 10956 15568 10968
rect 15620 10996 15626 11008
rect 16592 10996 16620 11036
rect 17129 11033 17141 11036
rect 17175 11033 17187 11067
rect 17129 11027 17187 11033
rect 15620 10968 16620 10996
rect 15620 10956 15626 10968
rect 552 10906 19412 10928
rect 552 10854 2755 10906
rect 2807 10854 2819 10906
rect 2871 10854 2883 10906
rect 2935 10854 2947 10906
rect 2999 10854 3011 10906
rect 3063 10854 7470 10906
rect 7522 10854 7534 10906
rect 7586 10854 7598 10906
rect 7650 10854 7662 10906
rect 7714 10854 7726 10906
rect 7778 10854 12185 10906
rect 12237 10854 12249 10906
rect 12301 10854 12313 10906
rect 12365 10854 12377 10906
rect 12429 10854 12441 10906
rect 12493 10854 16900 10906
rect 16952 10854 16964 10906
rect 17016 10854 17028 10906
rect 17080 10854 17092 10906
rect 17144 10854 17156 10906
rect 17208 10854 19412 10906
rect 552 10832 19412 10854
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3142 10792 3148 10804
rect 3099 10764 3148 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9548 10764 9781 10792
rect 9548 10752 9554 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 13262 10752 13268 10804
rect 13320 10792 13326 10804
rect 14093 10795 14151 10801
rect 14093 10792 14105 10795
rect 13320 10764 14105 10792
rect 13320 10752 13326 10764
rect 14093 10761 14105 10764
rect 14139 10761 14151 10795
rect 14093 10755 14151 10761
rect 14458 10752 14464 10804
rect 14516 10752 14522 10804
rect 14734 10752 14740 10804
rect 14792 10792 14798 10804
rect 15470 10792 15476 10804
rect 14792 10764 15476 10792
rect 14792 10752 14798 10764
rect 15470 10752 15476 10764
rect 15528 10792 15534 10804
rect 15838 10792 15844 10804
rect 15528 10764 15844 10792
rect 15528 10752 15534 10764
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 11238 10724 11244 10736
rect 9732 10696 11244 10724
rect 9732 10684 9738 10696
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 11793 10727 11851 10733
rect 11793 10693 11805 10727
rect 11839 10724 11851 10727
rect 13446 10724 13452 10736
rect 11839 10696 13452 10724
rect 11839 10693 11851 10696
rect 11793 10687 11851 10693
rect 12820 10668 12848 10696
rect 13446 10684 13452 10696
rect 13504 10684 13510 10736
rect 14182 10724 14188 10736
rect 13648 10696 14188 10724
rect 8018 10656 8024 10668
rect 7576 10628 8024 10656
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 1762 10588 1768 10600
rect 1719 10560 1768 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 1940 10591 1998 10597
rect 1940 10557 1952 10591
rect 1986 10557 1998 10591
rect 1940 10551 1998 10557
rect 1854 10480 1860 10532
rect 1912 10520 1918 10532
rect 1964 10520 1992 10551
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7576 10597 7604 10628
rect 8018 10616 8024 10628
rect 8076 10616 8082 10668
rect 11330 10616 11336 10668
rect 11388 10616 11394 10668
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 13648 10600 13676 10696
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 15010 10724 15016 10736
rect 14292 10696 15016 10724
rect 14292 10656 14320 10696
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15286 10724 15292 10736
rect 15120 10696 15292 10724
rect 15120 10656 15148 10696
rect 15286 10684 15292 10696
rect 15344 10684 15350 10736
rect 17129 10727 17187 10733
rect 16316 10696 16620 10724
rect 16316 10668 16344 10696
rect 14108 10628 14320 10656
rect 14752 10628 15148 10656
rect 14001 10601 14059 10607
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7432 10560 7573 10588
rect 7432 10548 7438 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 7926 10588 7932 10600
rect 7791 10560 7932 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8386 10548 8392 10600
rect 8444 10548 8450 10600
rect 8656 10591 8714 10597
rect 8656 10557 8668 10591
rect 8702 10588 8714 10591
rect 9030 10588 9036 10600
rect 8702 10560 9036 10588
rect 8702 10557 8714 10560
rect 8656 10551 8714 10557
rect 9030 10548 9036 10560
rect 9088 10548 9094 10600
rect 11422 10548 11428 10600
rect 11480 10588 11486 10600
rect 12618 10588 12624 10600
rect 11480 10560 12624 10588
rect 11480 10548 11486 10560
rect 12618 10548 12624 10560
rect 12676 10548 12682 10600
rect 13541 10591 13599 10597
rect 13541 10557 13553 10591
rect 13587 10588 13599 10591
rect 13630 10588 13636 10600
rect 13587 10560 13636 10588
rect 13587 10557 13599 10560
rect 13541 10551 13599 10557
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10557 13783 10591
rect 13725 10551 13783 10557
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10590 13875 10591
rect 13863 10562 13952 10590
rect 13863 10557 13875 10562
rect 13817 10551 13875 10557
rect 1912 10492 1992 10520
rect 1912 10480 1918 10492
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 13740 10520 13768 10551
rect 13412 10492 13768 10520
rect 13924 10520 13952 10562
rect 14001 10567 14013 10601
rect 14047 10598 14059 10601
rect 14108 10598 14136 10628
rect 14047 10570 14136 10598
rect 14047 10567 14059 10570
rect 14001 10561 14059 10567
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14240 10560 14289 10588
rect 14240 10548 14246 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14553 10591 14611 10597
rect 14553 10557 14565 10591
rect 14599 10588 14611 10591
rect 14752 10588 14780 10628
rect 15654 10616 15660 10668
rect 15712 10656 15718 10668
rect 16298 10656 16304 10668
rect 15712 10628 16304 10656
rect 15712 10616 15718 10628
rect 14599 10560 14780 10588
rect 14829 10591 14887 10597
rect 14599 10557 14611 10560
rect 14553 10551 14611 10557
rect 14829 10557 14841 10591
rect 14875 10557 14887 10591
rect 14829 10551 14887 10557
rect 14844 10520 14872 10551
rect 14918 10548 14924 10600
rect 14976 10548 14982 10600
rect 15013 10591 15071 10597
rect 15013 10557 15025 10591
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 13924 10492 14872 10520
rect 15028 10520 15056 10551
rect 15102 10548 15108 10600
rect 15160 10548 15166 10600
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10588 15807 10591
rect 15838 10588 15844 10600
rect 15795 10560 15844 10588
rect 15795 10557 15807 10560
rect 15749 10551 15807 10557
rect 15838 10548 15844 10560
rect 15896 10548 15902 10600
rect 15948 10597 15976 10628
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16592 10665 16620 10696
rect 17129 10693 17141 10727
rect 17175 10724 17187 10727
rect 17218 10724 17224 10736
rect 17175 10696 17224 10724
rect 17175 10693 17187 10696
rect 17129 10687 17187 10693
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 16485 10659 16543 10665
rect 16485 10656 16497 10659
rect 16448 10628 16497 10656
rect 16448 10616 16454 10628
rect 16485 10625 16497 10628
rect 16531 10625 16543 10659
rect 16485 10619 16543 10625
rect 16577 10659 16635 10665
rect 16577 10625 16589 10659
rect 16623 10625 16635 10659
rect 16577 10619 16635 10625
rect 15933 10591 15991 10597
rect 15933 10557 15945 10591
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16816 10560 16957 10588
rect 16816 10548 16822 10560
rect 16945 10557 16957 10560
rect 16991 10588 17003 10591
rect 17494 10588 17500 10600
rect 16991 10560 17500 10588
rect 16991 10557 17003 10560
rect 16945 10551 17003 10557
rect 17494 10548 17500 10560
rect 17552 10548 17558 10600
rect 15028 10492 15148 10520
rect 13412 10480 13418 10492
rect 14016 10464 14044 10492
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 8294 10452 8300 10464
rect 7791 10424 8300 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8294 10412 8300 10424
rect 8352 10412 8358 10464
rect 13538 10412 13544 10464
rect 13596 10412 13602 10464
rect 13906 10412 13912 10464
rect 13964 10412 13970 10464
rect 13998 10412 14004 10464
rect 14056 10412 14062 10464
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 14424 10424 14657 10452
rect 14424 10412 14430 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 14844 10452 14872 10492
rect 15010 10452 15016 10464
rect 14844 10424 15016 10452
rect 14645 10415 14703 10421
rect 15010 10412 15016 10424
rect 15068 10412 15074 10464
rect 15120 10452 15148 10492
rect 15194 10452 15200 10464
rect 15120 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10452 15258 10464
rect 15838 10452 15844 10464
rect 15252 10424 15844 10452
rect 15252 10412 15258 10424
rect 15838 10412 15844 10424
rect 15896 10412 15902 10464
rect 16022 10412 16028 10464
rect 16080 10412 16086 10464
rect 16393 10455 16451 10461
rect 16393 10421 16405 10455
rect 16439 10452 16451 10455
rect 16482 10452 16488 10464
rect 16439 10424 16488 10452
rect 16439 10421 16451 10424
rect 16393 10415 16451 10421
rect 16482 10412 16488 10424
rect 16540 10452 16546 10464
rect 17862 10452 17868 10464
rect 16540 10424 17868 10452
rect 16540 10412 16546 10424
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 552 10362 19571 10384
rect 552 10310 5112 10362
rect 5164 10310 5176 10362
rect 5228 10310 5240 10362
rect 5292 10310 5304 10362
rect 5356 10310 5368 10362
rect 5420 10310 9827 10362
rect 9879 10310 9891 10362
rect 9943 10310 9955 10362
rect 10007 10310 10019 10362
rect 10071 10310 10083 10362
rect 10135 10310 14542 10362
rect 14594 10310 14606 10362
rect 14658 10310 14670 10362
rect 14722 10310 14734 10362
rect 14786 10310 14798 10362
rect 14850 10310 19257 10362
rect 19309 10310 19321 10362
rect 19373 10310 19385 10362
rect 19437 10310 19449 10362
rect 19501 10310 19513 10362
rect 19565 10310 19571 10362
rect 552 10288 19571 10310
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 10686 10248 10692 10260
rect 7055 10220 10692 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 13630 10208 13636 10260
rect 13688 10208 13694 10260
rect 14182 10208 14188 10260
rect 14240 10208 14246 10260
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 15194 10248 15200 10260
rect 14323 10220 15200 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 15378 10208 15384 10260
rect 15436 10248 15442 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 15436 10220 17785 10248
rect 15436 10208 15442 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 17862 10208 17868 10260
rect 17920 10208 17926 10260
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 9876 10152 10425 10180
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7006 10112 7012 10124
rect 6963 10084 7012 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7374 10112 7380 10124
rect 7147 10084 7380 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 7561 10115 7619 10121
rect 7561 10081 7573 10115
rect 7607 10112 7619 10115
rect 8202 10112 8208 10124
rect 7607 10084 8208 10112
rect 7607 10081 7619 10084
rect 7561 10075 7619 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9876 10121 9904 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 13648 10180 13676 10208
rect 10413 10143 10471 10149
rect 13372 10152 13676 10180
rect 9861 10115 9919 10121
rect 9861 10112 9873 10115
rect 9548 10084 9873 10112
rect 9548 10072 9554 10084
rect 9861 10081 9873 10084
rect 9907 10081 9919 10115
rect 9861 10075 9919 10081
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 10008 10084 10057 10112
rect 10008 10072 10014 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10192 10084 10241 10112
rect 10192 10072 10198 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 10229 10075 10287 10081
rect 11238 10072 11244 10124
rect 11296 10072 11302 10124
rect 11977 10115 12035 10121
rect 11977 10081 11989 10115
rect 12023 10112 12035 10115
rect 12618 10112 12624 10124
rect 12023 10084 12624 10112
rect 12023 10081 12035 10084
rect 11977 10075 12035 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 13262 10072 13268 10124
rect 13320 10072 13326 10124
rect 13372 10121 13400 10152
rect 13906 10140 13912 10192
rect 13964 10180 13970 10192
rect 14553 10183 14611 10189
rect 14553 10180 14565 10183
rect 13964 10152 14565 10180
rect 13964 10140 13970 10152
rect 14553 10149 14565 10152
rect 14599 10149 14611 10183
rect 14553 10143 14611 10149
rect 15746 10140 15752 10192
rect 15804 10180 15810 10192
rect 16022 10180 16028 10192
rect 15804 10152 16028 10180
rect 15804 10140 15810 10152
rect 16022 10140 16028 10152
rect 16080 10180 16086 10192
rect 16117 10183 16175 10189
rect 16117 10180 16129 10183
rect 16080 10152 16129 10180
rect 16080 10140 16086 10152
rect 16117 10149 16129 10152
rect 16163 10149 16175 10183
rect 16117 10143 16175 10149
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10081 13415 10115
rect 13357 10075 13415 10081
rect 13630 10072 13636 10124
rect 13688 10072 13694 10124
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10081 14519 10115
rect 14461 10075 14519 10081
rect 7392 9976 7420 10072
rect 9766 10004 9772 10056
rect 9824 10044 9830 10056
rect 10318 10044 10324 10056
rect 9824 10016 10324 10044
rect 9824 10004 9830 10016
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10044 13507 10047
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13495 10016 13737 10044
rect 13495 10013 13507 10016
rect 13449 10007 13507 10013
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 10134 9976 10140 9988
rect 7392 9948 10140 9976
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 12894 9936 12900 9988
rect 12952 9976 12958 9988
rect 13924 9976 13952 10007
rect 13998 10004 14004 10056
rect 14056 10004 14062 10056
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14476 10044 14504 10075
rect 14642 10072 14648 10124
rect 14700 10112 14706 10124
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14700 10084 14749 10112
rect 14700 10072 14706 10084
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 14752 10044 14780 10075
rect 16206 10072 16212 10124
rect 16264 10112 16270 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 16264 10084 16313 10112
rect 16264 10072 16270 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10112 16451 10115
rect 17310 10112 17316 10124
rect 16439 10084 17316 10112
rect 16439 10081 16451 10084
rect 16393 10075 16451 10081
rect 17310 10072 17316 10084
rect 17368 10072 17374 10124
rect 16114 10044 16120 10056
rect 14476 10016 14596 10044
rect 14752 10016 16120 10044
rect 12952 9948 13952 9976
rect 12952 9936 12958 9948
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7469 9911 7527 9917
rect 7469 9908 7481 9911
rect 7432 9880 7481 9908
rect 7432 9868 7438 9880
rect 7469 9877 7481 9880
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 10505 9911 10563 9917
rect 10505 9908 10517 9911
rect 9548 9880 10517 9908
rect 9548 9868 9554 9880
rect 10505 9877 10517 9880
rect 10551 9877 10563 9911
rect 10505 9871 10563 9877
rect 12986 9868 12992 9920
rect 13044 9868 13050 9920
rect 13262 9868 13268 9920
rect 13320 9908 13326 9920
rect 14568 9908 14596 10016
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 14734 9936 14740 9988
rect 14792 9936 14798 9988
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 17972 9976 18000 10007
rect 16632 9948 18000 9976
rect 16632 9936 16638 9948
rect 17880 9920 17908 9948
rect 13320 9880 14596 9908
rect 16117 9911 16175 9917
rect 13320 9868 13326 9880
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16298 9908 16304 9920
rect 16163 9880 16304 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 17310 9868 17316 9920
rect 17368 9908 17374 9920
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17368 9880 17417 9908
rect 17368 9868 17374 9880
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17405 9871 17463 9877
rect 17862 9868 17868 9920
rect 17920 9868 17926 9920
rect 552 9818 19412 9840
rect 552 9766 2755 9818
rect 2807 9766 2819 9818
rect 2871 9766 2883 9818
rect 2935 9766 2947 9818
rect 2999 9766 3011 9818
rect 3063 9766 7470 9818
rect 7522 9766 7534 9818
rect 7586 9766 7598 9818
rect 7650 9766 7662 9818
rect 7714 9766 7726 9818
rect 7778 9766 12185 9818
rect 12237 9766 12249 9818
rect 12301 9766 12313 9818
rect 12365 9766 12377 9818
rect 12429 9766 12441 9818
rect 12493 9766 16900 9818
rect 16952 9766 16964 9818
rect 17016 9766 17028 9818
rect 17080 9766 17092 9818
rect 17144 9766 17156 9818
rect 17208 9766 19412 9818
rect 552 9744 19412 9766
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10226 9704 10232 9716
rect 10008 9676 10232 9704
rect 10008 9664 10014 9676
rect 10226 9664 10232 9676
rect 10284 9704 10290 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 10284 9676 10517 9704
rect 10284 9664 10290 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 10505 9667 10563 9673
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 13817 9707 13875 9713
rect 13817 9704 13829 9707
rect 12676 9676 13829 9704
rect 12676 9664 12682 9676
rect 13817 9673 13829 9676
rect 13863 9673 13875 9707
rect 13817 9667 13875 9673
rect 12986 9636 12992 9648
rect 9140 9608 12992 9636
rect 7929 9571 7987 9577
rect 7929 9537 7941 9571
rect 7975 9568 7987 9571
rect 8386 9568 8392 9580
rect 7975 9540 8392 9568
rect 7975 9537 7987 9540
rect 7929 9531 7987 9537
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 9140 9577 9168 9608
rect 12986 9596 12992 9608
rect 13044 9596 13050 9648
rect 13832 9636 13860 9667
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 14366 9704 14372 9716
rect 14148 9676 14372 9704
rect 14148 9664 14154 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 14476 9676 15148 9704
rect 14476 9636 14504 9676
rect 13832 9608 14504 9636
rect 15120 9636 15148 9676
rect 15194 9664 15200 9716
rect 15252 9704 15258 9716
rect 16482 9704 16488 9716
rect 15252 9676 16488 9704
rect 15252 9664 15258 9676
rect 16482 9664 16488 9676
rect 16540 9664 16546 9716
rect 16666 9636 16672 9648
rect 15120 9608 16672 9636
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 9125 9571 9183 9577
rect 9125 9537 9137 9571
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 11057 9571 11115 9577
rect 10367 9540 10916 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 8987 9472 9689 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9677 9469 9689 9472
rect 9723 9500 9735 9503
rect 9766 9500 9772 9512
rect 9723 9472 9772 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 7650 9392 7656 9444
rect 7708 9441 7714 9444
rect 7708 9395 7720 9441
rect 7708 9392 7714 9395
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6236 9336 6561 9364
rect 6236 9324 6242 9336
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6549 9327 6607 9333
rect 7466 9324 7472 9376
rect 7524 9364 7530 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 7524 9336 8493 9364
rect 7524 9324 7530 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9490 9364 9496 9376
rect 8895 9336 9496 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9876 9364 9904 9463
rect 9950 9460 9956 9512
rect 10008 9460 10014 9512
rect 10042 9460 10048 9512
rect 10100 9460 10106 9512
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 10405 9503 10463 9509
rect 10405 9500 10417 9503
rect 10192 9472 10417 9500
rect 10192 9460 10198 9472
rect 10405 9469 10417 9472
rect 10451 9469 10463 9503
rect 10405 9463 10463 9469
rect 10888 9432 10916 9540
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11422 9568 11428 9580
rect 11103 9540 11428 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 11422 9528 11428 9540
rect 11480 9528 11486 9580
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12710 9568 12716 9580
rect 11931 9540 12716 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12710 9528 12716 9540
rect 12768 9568 12774 9580
rect 13170 9568 13176 9580
rect 12768 9540 13176 9568
rect 12768 9528 12774 9540
rect 13170 9528 13176 9540
rect 13228 9528 13234 9580
rect 14458 9568 14464 9580
rect 14108 9540 14464 9568
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 12406 9472 13676 9500
rect 12406 9432 12434 9472
rect 10888 9404 12434 9432
rect 10410 9364 10416 9376
rect 9876 9336 10416 9364
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 11940 9336 13553 9364
rect 11940 9324 11946 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 13648 9364 13676 9472
rect 13722 9460 13728 9512
rect 13780 9460 13786 9512
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14108 9500 14136 9540
rect 14458 9528 14464 9540
rect 14516 9568 14522 9580
rect 15378 9568 15384 9580
rect 14516 9540 15384 9568
rect 14516 9528 14522 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 17310 9568 17316 9580
rect 16224 9540 17316 9568
rect 14047 9472 14136 9500
rect 14185 9503 14243 9509
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 15194 9500 15200 9512
rect 14231 9472 15200 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 15746 9460 15752 9512
rect 15804 9500 15810 9512
rect 15933 9503 15991 9509
rect 15933 9500 15945 9503
rect 15804 9472 15945 9500
rect 15804 9460 15810 9472
rect 15933 9469 15945 9472
rect 15979 9469 15991 9503
rect 15933 9463 15991 9469
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16224 9500 16252 9540
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 16071 9472 16252 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16298 9460 16304 9512
rect 16356 9460 16362 9512
rect 16393 9503 16451 9509
rect 16393 9469 16405 9503
rect 16439 9500 16451 9503
rect 16666 9500 16672 9512
rect 16439 9472 16672 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 13740 9432 13768 9460
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 13740 9404 16129 9432
rect 16117 9401 16129 9404
rect 16163 9432 16175 9435
rect 16206 9432 16212 9444
rect 16163 9404 16212 9432
rect 16163 9401 16175 9404
rect 16117 9395 16175 9401
rect 16206 9392 16212 9404
rect 16264 9392 16270 9444
rect 15194 9364 15200 9376
rect 13648 9336 15200 9364
rect 13541 9327 13599 9333
rect 15194 9324 15200 9336
rect 15252 9324 15258 9376
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15749 9367 15807 9373
rect 15749 9364 15761 9367
rect 15344 9336 15761 9364
rect 15344 9324 15350 9336
rect 15749 9333 15761 9336
rect 15795 9333 15807 9367
rect 15749 9327 15807 9333
rect 552 9274 19571 9296
rect 552 9222 5112 9274
rect 5164 9222 5176 9274
rect 5228 9222 5240 9274
rect 5292 9222 5304 9274
rect 5356 9222 5368 9274
rect 5420 9222 9827 9274
rect 9879 9222 9891 9274
rect 9943 9222 9955 9274
rect 10007 9222 10019 9274
rect 10071 9222 10083 9274
rect 10135 9222 14542 9274
rect 14594 9222 14606 9274
rect 14658 9222 14670 9274
rect 14722 9222 14734 9274
rect 14786 9222 14798 9274
rect 14850 9222 19257 9274
rect 19309 9222 19321 9274
rect 19373 9222 19385 9274
rect 19437 9222 19449 9274
rect 19501 9222 19513 9274
rect 19565 9222 19571 9274
rect 552 9200 19571 9222
rect 7374 9120 7380 9172
rect 7432 9160 7438 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 7432 9132 7481 9160
rect 7432 9120 7438 9132
rect 7469 9129 7481 9132
rect 7515 9129 7527 9163
rect 7469 9123 7527 9129
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 10229 9163 10287 9169
rect 10229 9160 10241 9163
rect 9079 9132 10241 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 10229 9129 10241 9132
rect 10275 9129 10287 9163
rect 10229 9123 10287 9129
rect 11514 9120 11520 9172
rect 11572 9160 11578 9172
rect 12894 9160 12900 9172
rect 11572 9132 12900 9160
rect 11572 9120 11578 9132
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 13262 9120 13268 9172
rect 13320 9120 13326 9172
rect 15841 9163 15899 9169
rect 15841 9129 15853 9163
rect 15887 9160 15899 9163
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 15887 9132 16129 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16117 9129 16129 9132
rect 16163 9129 16175 9163
rect 16117 9123 16175 9129
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 7653 9095 7711 9101
rect 7653 9061 7665 9095
rect 7699 9092 7711 9095
rect 8849 9095 8907 9101
rect 8849 9092 8861 9095
rect 7699 9064 8861 9092
rect 7699 9061 7711 9064
rect 7653 9055 7711 9061
rect 8849 9061 8861 9064
rect 8895 9092 8907 9095
rect 8938 9092 8944 9104
rect 8895 9064 8944 9092
rect 8895 9061 8907 9064
rect 8849 9055 8907 9061
rect 8938 9052 8944 9064
rect 8996 9052 9002 9104
rect 11977 9095 12035 9101
rect 11977 9092 11989 9095
rect 9692 9064 11989 9092
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 9024 7435 9027
rect 7466 9024 7472 9036
rect 7423 8996 7472 9024
rect 7423 8993 7435 8996
rect 7377 8987 7435 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 9171 8996 9352 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 9324 8965 9352 8996
rect 9490 8984 9496 9036
rect 9548 8984 9554 9036
rect 9692 9033 9720 9064
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10226 9024 10232 9036
rect 9999 8996 10232 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10336 9033 10364 9064
rect 11977 9061 11989 9064
rect 12023 9061 12035 9095
rect 11977 9055 12035 9061
rect 12437 9095 12495 9101
rect 12437 9061 12449 9095
rect 12483 9092 12495 9095
rect 16960 9092 16988 9123
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17313 9163 17371 9169
rect 17313 9160 17325 9163
rect 17276 9132 17325 9160
rect 17276 9120 17282 9132
rect 17313 9129 17325 9132
rect 17359 9129 17371 9163
rect 17313 9123 17371 9129
rect 12483 9064 16988 9092
rect 17957 9095 18015 9101
rect 12483 9061 12495 9064
rect 12437 9055 12495 9061
rect 17957 9061 17969 9095
rect 18003 9061 18015 9095
rect 17957 9055 18015 9061
rect 10321 9027 10379 9033
rect 10321 8993 10333 9027
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 9309 8959 9367 8965
rect 9309 8925 9321 8959
rect 9355 8925 9367 8959
rect 9309 8919 9367 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 10410 8956 10416 8968
rect 9815 8928 10416 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10520 8956 10548 8987
rect 11514 8984 11520 9036
rect 11572 9024 11578 9036
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11572 8996 11621 9024
rect 11572 8984 11578 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11790 8984 11796 9036
rect 11848 8984 11854 9036
rect 11882 8984 11888 9036
rect 11940 8984 11946 9036
rect 12253 9027 12311 9033
rect 12253 9024 12265 9027
rect 11992 8996 12265 9024
rect 10520 8928 11652 8956
rect 7650 8848 7656 8900
rect 7708 8848 7714 8900
rect 9585 8891 9643 8897
rect 9585 8857 9597 8891
rect 9631 8888 9643 8891
rect 10520 8888 10548 8928
rect 11624 8897 11652 8928
rect 9631 8860 10548 8888
rect 11609 8891 11667 8897
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 11609 8857 11621 8891
rect 11655 8857 11667 8891
rect 11992 8888 12020 8996
rect 12253 8993 12265 8996
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 13078 9024 13084 9036
rect 12584 8996 13084 9024
rect 12584 8984 12590 8996
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 13170 8984 13176 9036
rect 13228 8984 13234 9036
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 13722 9024 13728 9036
rect 13587 8996 13728 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 15654 8984 15660 9036
rect 15712 8984 15718 9036
rect 15930 8984 15936 9036
rect 15988 8984 15994 9036
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 9024 16727 9027
rect 17310 9024 17316 9036
rect 16715 8996 17316 9024
rect 16715 8993 16727 8996
rect 16669 8987 16727 8993
rect 17310 8984 17316 8996
rect 17368 9024 17374 9036
rect 17972 9024 18000 9055
rect 17368 8996 18000 9024
rect 18141 9027 18199 9033
rect 17368 8984 17374 8996
rect 18141 8993 18153 9027
rect 18187 9024 18199 9027
rect 18322 9024 18328 9036
rect 18187 8996 18328 9024
rect 18187 8993 18199 8996
rect 18141 8987 18199 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 12069 8959 12127 8965
rect 12069 8925 12081 8959
rect 12115 8956 12127 8959
rect 12710 8956 12716 8968
rect 12115 8928 12716 8956
rect 12115 8925 12127 8928
rect 12069 8919 12127 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 15838 8956 15844 8968
rect 13495 8928 15844 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16393 8959 16451 8965
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 17218 8956 17224 8968
rect 16439 8928 17224 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 12618 8888 12624 8900
rect 11992 8860 12624 8888
rect 11609 8851 11667 8857
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 15010 8848 15016 8900
rect 15068 8888 15074 8900
rect 16408 8888 16436 8919
rect 17218 8916 17224 8928
rect 17276 8916 17282 8968
rect 17402 8916 17408 8968
rect 17460 8916 17466 8968
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 17635 8928 17785 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17773 8925 17785 8928
rect 17819 8925 17831 8959
rect 17773 8919 17831 8925
rect 15068 8860 16436 8888
rect 15068 8848 15074 8860
rect 8846 8780 8852 8832
rect 8904 8780 8910 8832
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10318 8820 10324 8832
rect 10091 8792 10324 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 12161 8823 12219 8829
rect 12161 8789 12173 8823
rect 12207 8820 12219 8823
rect 12805 8823 12863 8829
rect 12805 8820 12817 8823
rect 12207 8792 12817 8820
rect 12207 8789 12219 8792
rect 12161 8783 12219 8789
rect 12805 8789 12817 8792
rect 12851 8789 12863 8823
rect 12805 8783 12863 8789
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 15657 8823 15715 8829
rect 15657 8820 15669 8823
rect 15436 8792 15669 8820
rect 15436 8780 15442 8792
rect 15657 8789 15669 8792
rect 15703 8789 15715 8823
rect 15657 8783 15715 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16301 8823 16359 8829
rect 16301 8820 16313 8823
rect 16172 8792 16313 8820
rect 16172 8780 16178 8792
rect 16301 8789 16313 8792
rect 16347 8789 16359 8823
rect 16301 8783 16359 8789
rect 552 8730 19412 8752
rect 552 8678 2755 8730
rect 2807 8678 2819 8730
rect 2871 8678 2883 8730
rect 2935 8678 2947 8730
rect 2999 8678 3011 8730
rect 3063 8678 7470 8730
rect 7522 8678 7534 8730
rect 7586 8678 7598 8730
rect 7650 8678 7662 8730
rect 7714 8678 7726 8730
rect 7778 8678 12185 8730
rect 12237 8678 12249 8730
rect 12301 8678 12313 8730
rect 12365 8678 12377 8730
rect 12429 8678 12441 8730
rect 12493 8678 16900 8730
rect 16952 8678 16964 8730
rect 17016 8678 17028 8730
rect 17080 8678 17092 8730
rect 17144 8678 17156 8730
rect 17208 8678 19412 8730
rect 552 8656 19412 8678
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 11848 8588 12265 8616
rect 11848 8576 11854 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13228 8588 13277 8616
rect 13228 8576 13234 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 14090 8576 14096 8628
rect 14148 8616 14154 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 14148 8588 16313 8616
rect 14148 8576 14154 8588
rect 16301 8585 16313 8588
rect 16347 8616 16359 8619
rect 16758 8616 16764 8628
rect 16347 8588 16764 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 17405 8619 17463 8625
rect 17405 8585 17417 8619
rect 17451 8585 17463 8619
rect 18322 8616 18328 8628
rect 17405 8579 17463 8585
rect 17880 8588 18328 8616
rect 8481 8551 8539 8557
rect 8481 8517 8493 8551
rect 8527 8548 8539 8551
rect 8662 8548 8668 8560
rect 8527 8520 8668 8548
rect 8527 8517 8539 8520
rect 8481 8511 8539 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 15010 8548 15016 8560
rect 14108 8520 15016 8548
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13320 8452 13737 8480
rect 13320 8440 13326 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 8444 8384 9873 8412
rect 8444 8372 8450 8384
rect 9861 8381 9873 8384
rect 9907 8412 9919 8415
rect 11977 8415 12035 8421
rect 11977 8412 11989 8415
rect 9907 8384 11989 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 11977 8381 11989 8384
rect 12023 8381 12035 8415
rect 11977 8375 12035 8381
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 13170 8372 13176 8424
rect 13228 8372 13234 8424
rect 13357 8415 13415 8421
rect 13357 8381 13369 8415
rect 13403 8412 13415 8415
rect 13814 8412 13820 8424
rect 13403 8384 13820 8412
rect 13403 8381 13415 8384
rect 13357 8375 13415 8381
rect 13814 8372 13820 8384
rect 13872 8372 13878 8424
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14108 8412 14136 8520
rect 15010 8508 15016 8520
rect 15068 8508 15074 8560
rect 17420 8548 17448 8579
rect 15212 8520 17448 8548
rect 17497 8551 17555 8557
rect 14918 8480 14924 8492
rect 14660 8452 14924 8480
rect 13955 8384 14136 8412
rect 14185 8415 14243 8421
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 14185 8381 14197 8415
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 8846 8304 8852 8356
rect 8904 8344 8910 8356
rect 9594 8347 9652 8353
rect 9594 8344 9606 8347
rect 8904 8316 9606 8344
rect 8904 8304 8910 8316
rect 9594 8313 9606 8316
rect 9640 8313 9652 8347
rect 9594 8307 9652 8313
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10413 8347 10471 8353
rect 10413 8344 10425 8347
rect 9824 8316 10425 8344
rect 9824 8304 9830 8316
rect 10413 8313 10425 8316
rect 10459 8313 10471 8347
rect 10413 8307 10471 8313
rect 12621 8347 12679 8353
rect 12621 8313 12633 8347
rect 12667 8344 12679 8347
rect 14200 8344 14228 8375
rect 14458 8372 14464 8424
rect 14516 8372 14522 8424
rect 14660 8421 14688 8452
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15212 8489 15240 8520
rect 17497 8517 17509 8551
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 16666 8440 16672 8492
rect 16724 8480 16730 8492
rect 17402 8480 17408 8492
rect 16724 8452 16804 8480
rect 16724 8440 16730 8452
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 14737 8415 14795 8421
rect 14737 8381 14749 8415
rect 14783 8412 14795 8415
rect 15105 8415 15163 8421
rect 14783 8384 15056 8412
rect 14783 8381 14795 8384
rect 14737 8375 14795 8381
rect 14277 8347 14335 8353
rect 14277 8344 14289 8347
rect 12667 8316 14289 8344
rect 12667 8313 12679 8316
rect 12621 8307 12679 8313
rect 14277 8313 14289 8316
rect 14323 8313 14335 8347
rect 14277 8307 14335 8313
rect 14090 8236 14096 8288
rect 14148 8236 14154 8288
rect 14918 8236 14924 8288
rect 14976 8236 14982 8288
rect 15028 8276 15056 8384
rect 15105 8381 15117 8415
rect 15151 8381 15163 8415
rect 15105 8375 15163 8381
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15654 8412 15660 8424
rect 15335 8384 15660 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 15120 8344 15148 8375
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15746 8372 15752 8424
rect 15804 8372 15810 8424
rect 15838 8372 15844 8424
rect 15896 8372 15902 8424
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 16485 8415 16543 8421
rect 16485 8381 16497 8415
rect 16531 8412 16543 8415
rect 16574 8412 16580 8424
rect 16531 8384 16580 8412
rect 16531 8381 16543 8384
rect 16485 8375 16543 8381
rect 16574 8372 16580 8384
rect 16632 8372 16638 8424
rect 16776 8421 16804 8452
rect 16960 8452 17408 8480
rect 16761 8415 16819 8421
rect 16761 8381 16773 8415
rect 16807 8381 16819 8415
rect 16761 8375 16819 8381
rect 16850 8372 16856 8424
rect 16908 8421 16914 8424
rect 16960 8421 16988 8452
rect 17402 8440 17408 8452
rect 17460 8440 17466 8492
rect 16908 8415 16988 8421
rect 16908 8381 16921 8415
rect 16955 8384 16988 8415
rect 16955 8381 16967 8384
rect 16908 8375 16967 8381
rect 16908 8372 16914 8375
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17267 8415 17325 8421
rect 17267 8381 17279 8415
rect 17313 8412 17325 8415
rect 17512 8412 17540 8511
rect 17880 8421 17908 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 18012 8452 18061 8480
rect 18012 8440 18018 8452
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 17313 8384 17540 8412
rect 17865 8415 17923 8421
rect 17313 8381 17325 8384
rect 17267 8375 17325 8381
rect 17865 8381 17877 8415
rect 17911 8381 17923 8415
rect 18325 8415 18383 8421
rect 18325 8412 18337 8415
rect 17865 8375 17923 8381
rect 17972 8384 18337 8412
rect 15565 8347 15623 8353
rect 15565 8344 15577 8347
rect 15120 8316 15577 8344
rect 15565 8313 15577 8316
rect 15611 8313 15623 8347
rect 15856 8344 15884 8372
rect 16390 8344 16396 8356
rect 15856 8316 16396 8344
rect 15565 8307 15623 8313
rect 16390 8304 16396 8316
rect 16448 8304 16454 8356
rect 16669 8347 16727 8353
rect 16669 8313 16681 8347
rect 16715 8313 16727 8347
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 16669 8307 16727 8313
rect 16776 8316 17049 8344
rect 15470 8276 15476 8288
rect 15028 8248 15476 8276
rect 15470 8236 15476 8248
rect 15528 8276 15534 8288
rect 16298 8276 16304 8288
rect 15528 8248 16304 8276
rect 15528 8236 15534 8248
rect 16298 8236 16304 8248
rect 16356 8276 16362 8288
rect 16684 8276 16712 8307
rect 16776 8288 16804 8316
rect 17037 8313 17049 8316
rect 17083 8313 17095 8347
rect 17037 8307 17095 8313
rect 16356 8248 16712 8276
rect 16356 8236 16362 8248
rect 16758 8236 16764 8288
rect 16816 8236 16822 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 17972 8285 18000 8384
rect 18325 8381 18337 8384
rect 18371 8381 18383 8415
rect 18325 8375 18383 8381
rect 18509 8415 18567 8421
rect 18509 8381 18521 8415
rect 18555 8381 18567 8415
rect 18509 8375 18567 8381
rect 18046 8304 18052 8356
rect 18104 8344 18110 8356
rect 18524 8344 18552 8375
rect 18104 8316 18552 8344
rect 18104 8304 18110 8316
rect 17957 8279 18015 8285
rect 17957 8276 17969 8279
rect 17920 8248 17969 8276
rect 17920 8236 17926 8248
rect 17957 8245 17969 8248
rect 18003 8245 18015 8279
rect 17957 8239 18015 8245
rect 552 8186 19571 8208
rect 552 8134 5112 8186
rect 5164 8134 5176 8186
rect 5228 8134 5240 8186
rect 5292 8134 5304 8186
rect 5356 8134 5368 8186
rect 5420 8134 9827 8186
rect 9879 8134 9891 8186
rect 9943 8134 9955 8186
rect 10007 8134 10019 8186
rect 10071 8134 10083 8186
rect 10135 8134 14542 8186
rect 14594 8134 14606 8186
rect 14658 8134 14670 8186
rect 14722 8134 14734 8186
rect 14786 8134 14798 8186
rect 14850 8134 19257 8186
rect 19309 8134 19321 8186
rect 19373 8134 19385 8186
rect 19437 8134 19449 8186
rect 19501 8134 19513 8186
rect 19565 8134 19571 8186
rect 552 8112 19571 8134
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9858 8072 9864 8084
rect 8987 8044 9864 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9858 8032 9864 8044
rect 9916 8072 9922 8084
rect 10318 8072 10324 8084
rect 9916 8044 10324 8072
rect 9916 8032 9922 8044
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 12618 8032 12624 8084
rect 12676 8032 12682 8084
rect 12710 8032 12716 8084
rect 12768 8072 12774 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12768 8044 13001 8072
rect 12768 8032 12774 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13357 8075 13415 8081
rect 13357 8041 13369 8075
rect 13403 8072 13415 8075
rect 13538 8072 13544 8084
rect 13403 8044 13544 8072
rect 13403 8041 13415 8044
rect 13357 8035 13415 8041
rect 8849 8007 8907 8013
rect 8849 7973 8861 8007
rect 8895 8004 8907 8007
rect 9490 8004 9496 8016
rect 8895 7976 9496 8004
rect 8895 7973 8907 7976
rect 8849 7967 8907 7973
rect 9490 7964 9496 7976
rect 9548 7964 9554 8016
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 13372 8004 13400 8035
rect 13538 8032 13544 8044
rect 13596 8032 13602 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15746 8072 15752 8084
rect 15611 8044 15752 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 15988 8044 16129 8072
rect 15988 8032 15994 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 16298 8032 16304 8084
rect 16356 8072 16362 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16356 8044 16957 8072
rect 16356 8032 16362 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 15010 8004 15016 8016
rect 12584 7976 13400 8004
rect 14568 7976 15016 8004
rect 12584 7964 12590 7976
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7936 12495 7939
rect 12894 7936 12900 7948
rect 12483 7908 12900 7936
rect 12483 7905 12495 7908
rect 12437 7899 12495 7905
rect 12894 7896 12900 7908
rect 12952 7896 12958 7948
rect 13170 7896 13176 7948
rect 13228 7896 13234 7948
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 13538 7936 13544 7948
rect 13495 7908 13544 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 14568 7945 14596 7976
rect 15010 7964 15016 7976
rect 15068 8004 15074 8016
rect 15764 8004 15792 8032
rect 16761 8007 16819 8013
rect 16761 8004 16773 8007
rect 15068 7976 15700 8004
rect 15764 7976 16344 8004
rect 15068 7964 15074 7976
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7905 14611 7939
rect 14553 7899 14611 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 15470 7936 15476 7948
rect 14783 7908 15476 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 15672 7936 15700 7976
rect 16316 7945 16344 7976
rect 16500 7976 16773 8004
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 15672 7908 15761 7936
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 16301 7939 16359 7945
rect 16301 7905 16313 7939
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 16390 7896 16396 7948
rect 16448 7896 16454 7948
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 13188 7868 13216 7896
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 13188 7840 14657 7868
rect 9125 7831 9183 7837
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 9140 7800 9168 7831
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 14884 7840 15945 7868
rect 14884 7828 14890 7840
rect 15933 7837 15945 7840
rect 15979 7868 15991 7871
rect 16500 7868 16528 7976
rect 16761 7973 16773 7976
rect 16807 8004 16819 8007
rect 17494 8004 17500 8016
rect 16807 7976 17500 8004
rect 16807 7973 16819 7976
rect 16761 7967 16819 7973
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 16574 7896 16580 7948
rect 16632 7896 16638 7948
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 16669 7899 16727 7905
rect 16960 7908 17049 7936
rect 15979 7840 16528 7868
rect 16684 7868 16712 7899
rect 16684 7840 16804 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 14918 7800 14924 7812
rect 9140 7772 14924 7800
rect 14918 7760 14924 7772
rect 14976 7760 14982 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 16574 7800 16580 7812
rect 15252 7772 16580 7800
rect 15252 7760 15258 7772
rect 16574 7760 16580 7772
rect 16632 7760 16638 7812
rect 16776 7809 16804 7840
rect 16761 7803 16819 7809
rect 16761 7769 16773 7803
rect 16807 7800 16819 7803
rect 16850 7800 16856 7812
rect 16807 7772 16856 7800
rect 16807 7769 16819 7772
rect 16761 7763 16819 7769
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 12894 7692 12900 7744
rect 12952 7732 12958 7744
rect 15010 7732 15016 7744
rect 12952 7704 15016 7732
rect 12952 7692 12958 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 16960 7732 16988 7908
rect 17037 7905 17049 7908
rect 17083 7936 17095 7939
rect 17862 7936 17868 7948
rect 17083 7908 17868 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 15160 7704 16988 7732
rect 15160 7692 15166 7704
rect 552 7642 19412 7664
rect 552 7590 2755 7642
rect 2807 7590 2819 7642
rect 2871 7590 2883 7642
rect 2935 7590 2947 7642
rect 2999 7590 3011 7642
rect 3063 7590 7470 7642
rect 7522 7590 7534 7642
rect 7586 7590 7598 7642
rect 7650 7590 7662 7642
rect 7714 7590 7726 7642
rect 7778 7590 12185 7642
rect 12237 7590 12249 7642
rect 12301 7590 12313 7642
rect 12365 7590 12377 7642
rect 12429 7590 12441 7642
rect 12493 7590 16900 7642
rect 16952 7590 16964 7642
rect 17016 7590 17028 7642
rect 17080 7590 17092 7642
rect 17144 7590 17156 7642
rect 17208 7590 19412 7642
rect 552 7568 19412 7590
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14826 7528 14832 7540
rect 13964 7500 14832 7528
rect 13964 7488 13970 7500
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 15749 7531 15807 7537
rect 15749 7528 15761 7531
rect 15620 7500 15761 7528
rect 15620 7488 15626 7500
rect 15749 7497 15761 7500
rect 15795 7497 15807 7531
rect 15749 7491 15807 7497
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16816 7500 16865 7528
rect 16816 7488 16822 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 8386 7460 8392 7472
rect 8220 7432 8392 7460
rect 8220 7401 8248 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8665 7463 8723 7469
rect 8665 7429 8677 7463
rect 8711 7429 8723 7463
rect 11609 7463 11667 7469
rect 11609 7460 11621 7463
rect 8665 7423 8723 7429
rect 9692 7432 11621 7460
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8680 7392 8708 7423
rect 9692 7401 9720 7432
rect 11609 7429 11621 7432
rect 11655 7429 11667 7463
rect 11609 7423 11667 7429
rect 8205 7355 8263 7361
rect 8312 7364 8708 7392
rect 9677 7395 9735 7401
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7324 7987 7327
rect 8312 7324 8340 7364
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 10505 7395 10563 7401
rect 10505 7361 10517 7395
rect 10551 7392 10563 7395
rect 10551 7364 11468 7392
rect 10551 7361 10563 7364
rect 10505 7355 10563 7361
rect 7975 7296 8340 7324
rect 8389 7327 8447 7333
rect 7975 7293 7987 7296
rect 7929 7287 7987 7293
rect 8389 7293 8401 7327
rect 8435 7324 8447 7327
rect 8478 7324 8484 7336
rect 8435 7296 8484 7324
rect 8435 7293 8447 7296
rect 8389 7287 8447 7293
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7324 8723 7327
rect 8938 7324 8944 7336
rect 8711 7296 8944 7324
rect 8711 7293 8723 7296
rect 8665 7287 8723 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9548 7296 9781 7324
rect 9548 7284 9554 7296
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 6546 7216 6552 7268
rect 6604 7216 6610 7268
rect 9784 7256 9812 7287
rect 9858 7284 9864 7336
rect 9916 7324 9922 7336
rect 10689 7327 10747 7333
rect 10689 7324 10701 7327
rect 9916 7296 10701 7324
rect 9916 7284 9922 7296
rect 10689 7293 10701 7296
rect 10735 7293 10747 7327
rect 10689 7287 10747 7293
rect 10597 7259 10655 7265
rect 10597 7256 10609 7259
rect 9784 7228 10609 7256
rect 10597 7225 10609 7228
rect 10643 7225 10655 7259
rect 10597 7219 10655 7225
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8352 7160 8493 7188
rect 8352 7148 8358 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8481 7151 8539 7157
rect 10229 7191 10287 7197
rect 10229 7157 10241 7191
rect 10275 7188 10287 7191
rect 10318 7188 10324 7200
rect 10275 7160 10324 7188
rect 10275 7157 10287 7160
rect 10229 7151 10287 7157
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 11054 7148 11060 7200
rect 11112 7148 11118 7200
rect 11440 7188 11468 7364
rect 11514 7284 11520 7336
rect 11572 7284 11578 7336
rect 11624 7256 11652 7423
rect 12802 7420 12808 7472
rect 12860 7460 12866 7472
rect 13170 7460 13176 7472
rect 12860 7432 13176 7460
rect 12860 7420 12866 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 15013 7463 15071 7469
rect 15013 7460 15025 7463
rect 14332 7432 15025 7460
rect 14332 7420 14338 7432
rect 15013 7429 15025 7432
rect 15059 7429 15071 7463
rect 16482 7460 16488 7472
rect 15013 7423 15071 7429
rect 15304 7432 16488 7460
rect 11716 7364 13308 7392
rect 11716 7333 11744 7364
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 11790 7284 11796 7336
rect 11848 7284 11854 7336
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7293 12035 7327
rect 11977 7287 12035 7293
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7324 12495 7327
rect 12618 7324 12624 7336
rect 12483 7296 12624 7324
rect 12483 7293 12495 7296
rect 12437 7287 12495 7293
rect 11992 7256 12020 7287
rect 12618 7284 12624 7296
rect 12676 7284 12682 7336
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 12986 7324 12992 7336
rect 12768 7296 12992 7324
rect 12768 7284 12774 7296
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13078 7284 13084 7336
rect 13136 7284 13142 7336
rect 13170 7284 13176 7336
rect 13228 7284 13234 7336
rect 11624 7228 12020 7256
rect 12066 7216 12072 7268
rect 12124 7216 12130 7268
rect 12158 7216 12164 7268
rect 12216 7216 12222 7268
rect 12299 7259 12357 7265
rect 12299 7225 12311 7259
rect 12345 7256 12357 7259
rect 12345 7228 12756 7256
rect 12345 7225 12357 7228
rect 12299 7219 12357 7225
rect 12529 7191 12587 7197
rect 12529 7188 12541 7191
rect 11440 7160 12541 7188
rect 12529 7157 12541 7160
rect 12575 7157 12587 7191
rect 12728 7188 12756 7228
rect 12802 7216 12808 7268
rect 12860 7216 12866 7268
rect 12897 7259 12955 7265
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 13280 7256 13308 7364
rect 13538 7352 13544 7404
rect 13596 7392 13602 7404
rect 13596 7364 14412 7392
rect 13596 7352 13602 7364
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 14001 7327 14059 7333
rect 13403 7296 13768 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 13446 7256 13452 7268
rect 12943 7228 13452 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 13740 7265 13768 7296
rect 14001 7293 14013 7327
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7225 13783 7259
rect 14016 7256 14044 7287
rect 14090 7284 14096 7336
rect 14148 7284 14154 7336
rect 14384 7333 14412 7364
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 15102 7392 15108 7404
rect 14516 7364 15108 7392
rect 14516 7352 14522 7364
rect 14185 7327 14243 7333
rect 14185 7293 14197 7327
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7293 14427 7327
rect 14369 7287 14427 7293
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 14826 7324 14832 7336
rect 14691 7296 14832 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14200 7256 14228 7287
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 14936 7333 14964 7364
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 15010 7284 15016 7336
rect 15068 7284 15074 7336
rect 15304 7333 15332 7432
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 16945 7395 17003 7401
rect 15611 7364 16712 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 16684 7336 16712 7364
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17218 7392 17224 7404
rect 16991 7364 17224 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 15120 7296 15301 7324
rect 14016 7228 14136 7256
rect 14200 7228 14504 7256
rect 13725 7219 13783 7225
rect 14108 7200 14136 7228
rect 14476 7200 14504 7228
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12728 7160 13277 7188
rect 12529 7151 12587 7157
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 14090 7148 14096 7200
rect 14148 7188 14154 7200
rect 14366 7188 14372 7200
rect 14148 7160 14372 7188
rect 14148 7148 14154 7160
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14458 7148 14464 7200
rect 14516 7148 14522 7200
rect 14829 7191 14887 7197
rect 14829 7157 14841 7191
rect 14875 7188 14887 7191
rect 15120 7188 15148 7296
rect 15289 7293 15301 7296
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 15838 7284 15844 7336
rect 15896 7284 15902 7336
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 15197 7259 15255 7265
rect 15197 7225 15209 7259
rect 15243 7256 15255 7259
rect 16960 7256 16988 7355
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 15243 7228 16988 7256
rect 15243 7225 15255 7228
rect 15197 7219 15255 7225
rect 14875 7160 15148 7188
rect 14875 7157 14887 7160
rect 14829 7151 14887 7157
rect 15562 7148 15568 7200
rect 15620 7148 15626 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 16485 7191 16543 7197
rect 16485 7188 16497 7191
rect 16448 7160 16497 7188
rect 16448 7148 16454 7160
rect 16485 7157 16497 7160
rect 16531 7157 16543 7191
rect 16485 7151 16543 7157
rect 552 7098 19571 7120
rect 552 7046 5112 7098
rect 5164 7046 5176 7098
rect 5228 7046 5240 7098
rect 5292 7046 5304 7098
rect 5356 7046 5368 7098
rect 5420 7046 9827 7098
rect 9879 7046 9891 7098
rect 9943 7046 9955 7098
rect 10007 7046 10019 7098
rect 10071 7046 10083 7098
rect 10135 7046 14542 7098
rect 14594 7046 14606 7098
rect 14658 7046 14670 7098
rect 14722 7046 14734 7098
rect 14786 7046 14798 7098
rect 14850 7046 19257 7098
rect 19309 7046 19321 7098
rect 19373 7046 19385 7098
rect 19437 7046 19449 7098
rect 19501 7046 19513 7098
rect 19565 7046 19571 7098
rect 552 7024 19571 7046
rect 9217 6987 9275 6993
rect 9217 6953 9229 6987
rect 9263 6984 9275 6987
rect 9674 6984 9680 6996
rect 9263 6956 9680 6984
rect 9263 6953 9275 6956
rect 9217 6947 9275 6953
rect 9674 6944 9680 6956
rect 9732 6984 9738 6996
rect 10321 6987 10379 6993
rect 10321 6984 10333 6987
rect 9732 6956 10333 6984
rect 9732 6944 9738 6956
rect 10321 6953 10333 6956
rect 10367 6953 10379 6987
rect 10321 6947 10379 6953
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 12124 6956 12265 6984
rect 12124 6944 12130 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 12618 6944 12624 6996
rect 12676 6944 12682 6996
rect 12897 6987 12955 6993
rect 12897 6953 12909 6987
rect 12943 6984 12955 6987
rect 13078 6984 13084 6996
rect 12943 6956 13084 6984
rect 12943 6953 12955 6956
rect 12897 6947 12955 6953
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13504 6956 13553 6984
rect 13504 6944 13510 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14274 6984 14280 6996
rect 13872 6956 14280 6984
rect 13872 6944 13878 6956
rect 14274 6944 14280 6956
rect 14332 6944 14338 6996
rect 8481 6919 8539 6925
rect 8481 6885 8493 6919
rect 8527 6916 8539 6919
rect 8938 6916 8944 6928
rect 8527 6888 8944 6916
rect 8527 6885 8539 6888
rect 8481 6879 8539 6885
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 9309 6919 9367 6925
rect 9309 6885 9321 6919
rect 9355 6916 9367 6919
rect 9490 6916 9496 6928
rect 9355 6888 9496 6916
rect 9355 6885 9367 6888
rect 9309 6879 9367 6885
rect 9490 6876 9496 6888
rect 9548 6916 9554 6928
rect 10229 6919 10287 6925
rect 10229 6916 10241 6919
rect 9548 6888 10241 6916
rect 9548 6876 9554 6888
rect 10229 6885 10241 6888
rect 10275 6885 10287 6919
rect 10229 6879 10287 6885
rect 11514 6876 11520 6928
rect 11572 6916 11578 6928
rect 12636 6916 12664 6944
rect 15562 6925 15568 6928
rect 14001 6919 14059 6925
rect 14001 6916 14013 6919
rect 11572 6888 12480 6916
rect 12636 6888 12848 6916
rect 11572 6876 11578 6888
rect 8570 6808 8576 6860
rect 8628 6848 8634 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8628 6820 8677 6848
rect 8628 6808 8634 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 8803 6820 8892 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 8864 6721 8892 6820
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6848 11115 6851
rect 11146 6848 11152 6860
rect 11103 6820 11152 6848
rect 11103 6817 11115 6820
rect 11057 6811 11115 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11241 6851 11299 6857
rect 11241 6817 11253 6851
rect 11287 6848 11299 6851
rect 11330 6848 11336 6860
rect 11287 6820 11336 6848
rect 11287 6817 11299 6820
rect 11241 6811 11299 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 12452 6857 12480 6888
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 12526 6848 12532 6860
rect 12483 6820 12532 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 12526 6808 12532 6820
rect 12584 6808 12590 6860
rect 12710 6808 12716 6860
rect 12768 6808 12774 6860
rect 12820 6857 12848 6888
rect 13556 6888 14013 6916
rect 13556 6860 13584 6888
rect 14001 6885 14013 6888
rect 14047 6885 14059 6919
rect 15519 6919 15568 6925
rect 14001 6879 14059 6885
rect 15120 6888 15424 6916
rect 12805 6851 12863 6857
rect 12805 6817 12817 6851
rect 12851 6817 12863 6851
rect 12805 6811 12863 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6780 10563 6783
rect 11790 6780 11796 6792
rect 10551 6752 11796 6780
rect 10551 6749 10563 6752
rect 10505 6743 10563 6749
rect 8849 6715 8907 6721
rect 8849 6681 8861 6715
rect 8895 6681 8907 6715
rect 9508 6712 9536 6743
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 13004 6780 13032 6811
rect 13538 6808 13544 6860
rect 13596 6808 13602 6860
rect 13725 6851 13783 6857
rect 13725 6817 13737 6851
rect 13771 6848 13783 6851
rect 13814 6848 13820 6860
rect 13771 6820 13820 6848
rect 13771 6817 13783 6820
rect 13725 6811 13783 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 13906 6808 13912 6860
rect 13964 6808 13970 6860
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 14274 6808 14280 6860
rect 14332 6808 14338 6860
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 14458 6848 14464 6860
rect 14415 6820 14464 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 14384 6780 14412 6811
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 14550 6808 14556 6860
rect 14608 6848 14614 6860
rect 15120 6848 15148 6888
rect 14608 6820 15148 6848
rect 14608 6808 14614 6820
rect 15194 6808 15200 6860
rect 15252 6808 15258 6860
rect 15286 6808 15292 6860
rect 15344 6808 15350 6860
rect 15396 6857 15424 6888
rect 15519 6885 15531 6919
rect 15565 6885 15568 6919
rect 15519 6879 15568 6885
rect 15562 6876 15568 6879
rect 15620 6876 15626 6928
rect 15654 6876 15660 6928
rect 15712 6876 15718 6928
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 15672 6848 15700 6876
rect 15427 6820 15700 6848
rect 16117 6851 16175 6857
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 16117 6817 16129 6851
rect 16163 6848 16175 6851
rect 16482 6848 16488 6860
rect 16163 6820 16488 6848
rect 16163 6817 16175 6820
rect 16117 6811 16175 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 13004 6752 14412 6780
rect 14568 6752 15669 6780
rect 14568 6721 14596 6752
rect 15657 6749 15669 6752
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16209 6783 16267 6789
rect 16209 6780 16221 6783
rect 16080 6752 16221 6780
rect 16080 6740 16086 6752
rect 16209 6749 16221 6752
rect 16255 6749 16267 6783
rect 16209 6743 16267 6749
rect 16390 6740 16396 6792
rect 16448 6740 16454 6792
rect 14553 6715 14611 6721
rect 9508 6684 14136 6712
rect 8849 6675 8907 6681
rect 8481 6647 8539 6653
rect 8481 6613 8493 6647
rect 8527 6644 8539 6647
rect 9582 6644 9588 6656
rect 8527 6616 9588 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 9950 6644 9956 6656
rect 9907 6616 9956 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 11238 6604 11244 6656
rect 11296 6604 11302 6656
rect 14108 6644 14136 6684
rect 14553 6681 14565 6715
rect 14599 6681 14611 6715
rect 14553 6675 14611 6681
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 16301 6715 16359 6721
rect 16301 6712 16313 6715
rect 15252 6684 16313 6712
rect 15252 6672 15258 6684
rect 16301 6681 16313 6684
rect 16347 6681 16359 6715
rect 16301 6675 16359 6681
rect 15013 6647 15071 6653
rect 15013 6644 15025 6647
rect 14108 6616 15025 6644
rect 15013 6613 15025 6616
rect 15059 6613 15071 6647
rect 15013 6607 15071 6613
rect 552 6554 19412 6576
rect 552 6502 2755 6554
rect 2807 6502 2819 6554
rect 2871 6502 2883 6554
rect 2935 6502 2947 6554
rect 2999 6502 3011 6554
rect 3063 6502 7470 6554
rect 7522 6502 7534 6554
rect 7586 6502 7598 6554
rect 7650 6502 7662 6554
rect 7714 6502 7726 6554
rect 7778 6502 12185 6554
rect 12237 6502 12249 6554
rect 12301 6502 12313 6554
rect 12365 6502 12377 6554
rect 12429 6502 12441 6554
rect 12493 6502 16900 6554
rect 16952 6502 16964 6554
rect 17016 6502 17028 6554
rect 17080 6502 17092 6554
rect 17144 6502 17156 6554
rect 17208 6502 19412 6554
rect 552 6480 19412 6502
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 8996 6412 10088 6440
rect 8996 6400 9002 6412
rect 8386 6196 8392 6248
rect 8444 6236 8450 6248
rect 9306 6236 9312 6248
rect 8444 6208 9312 6236
rect 8444 6196 8450 6208
rect 9306 6196 9312 6208
rect 9364 6236 9370 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9364 6208 9873 6236
rect 9364 6196 9370 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 9950 6196 9956 6248
rect 10008 6196 10014 6248
rect 10060 6236 10088 6412
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 14550 6440 14556 6452
rect 12584 6412 14556 6440
rect 12584 6400 12590 6412
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 10226 6332 10232 6384
rect 10284 6332 10290 6384
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11514 6372 11520 6384
rect 10643 6344 11520 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10060 6208 10241 6236
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 9582 6128 9588 6180
rect 9640 6177 9646 6180
rect 9640 6168 9652 6177
rect 10244 6168 10272 6199
rect 10318 6196 10324 6248
rect 10376 6196 10382 6248
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6236 10471 6239
rect 10686 6236 10692 6248
rect 10459 6208 10692 6236
rect 10459 6205 10471 6208
rect 10413 6199 10471 6205
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10597 6171 10655 6177
rect 10597 6168 10609 6171
rect 9640 6140 9685 6168
rect 10244 6140 10609 6168
rect 9640 6131 9652 6140
rect 10597 6137 10609 6140
rect 10643 6168 10655 6171
rect 11330 6168 11336 6180
rect 10643 6140 11336 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 9640 6128 9646 6131
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 8478 6060 8484 6112
rect 8536 6060 8542 6112
rect 9398 6060 9404 6112
rect 9456 6100 9462 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9456 6072 10057 6100
rect 9456 6060 9462 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 552 6010 19571 6032
rect 552 5958 5112 6010
rect 5164 5958 5176 6010
rect 5228 5958 5240 6010
rect 5292 5958 5304 6010
rect 5356 5958 5368 6010
rect 5420 5958 9827 6010
rect 9879 5958 9891 6010
rect 9943 5958 9955 6010
rect 10007 5958 10019 6010
rect 10071 5958 10083 6010
rect 10135 5958 14542 6010
rect 14594 5958 14606 6010
rect 14658 5958 14670 6010
rect 14722 5958 14734 6010
rect 14786 5958 14798 6010
rect 14850 5958 19257 6010
rect 19309 5958 19321 6010
rect 19373 5958 19385 6010
rect 19437 5958 19449 6010
rect 19501 5958 19513 6010
rect 19565 5958 19571 6010
rect 552 5936 19571 5958
rect 9324 5800 12434 5828
rect 9324 5772 9352 5800
rect 9306 5720 9312 5772
rect 9364 5720 9370 5772
rect 9576 5763 9634 5769
rect 9576 5729 9588 5763
rect 9622 5760 9634 5763
rect 10134 5760 10140 5772
rect 9622 5732 10140 5760
rect 9622 5729 9634 5732
rect 9576 5723 9634 5729
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 10980 5769 11008 5800
rect 10965 5763 11023 5769
rect 10965 5729 10977 5763
rect 11011 5760 11023 5763
rect 11054 5760 11060 5772
rect 11011 5732 11060 5760
rect 11011 5729 11023 5732
rect 10965 5723 11023 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11232 5763 11290 5769
rect 11232 5729 11244 5763
rect 11278 5760 11290 5763
rect 11514 5760 11520 5772
rect 11278 5732 11520 5760
rect 11278 5729 11290 5732
rect 11232 5723 11290 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 12406 5760 12434 5800
rect 16574 5788 16580 5840
rect 16632 5828 16638 5840
rect 17028 5831 17086 5837
rect 17028 5828 17040 5831
rect 16632 5800 17040 5828
rect 16632 5788 16638 5800
rect 17028 5797 17040 5800
rect 17074 5797 17086 5831
rect 17028 5791 17086 5797
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 12406 5732 16773 5760
rect 16761 5729 16773 5732
rect 16807 5729 16819 5763
rect 16761 5723 16819 5729
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5556 10747 5559
rect 11146 5556 11152 5568
rect 10735 5528 11152 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 12345 5559 12403 5565
rect 12345 5525 12357 5559
rect 12391 5556 12403 5559
rect 16114 5556 16120 5568
rect 12391 5528 16120 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 18141 5559 18199 5565
rect 18141 5525 18153 5559
rect 18187 5556 18199 5559
rect 18598 5556 18604 5568
rect 18187 5528 18604 5556
rect 18187 5525 18199 5528
rect 18141 5519 18199 5525
rect 18598 5516 18604 5528
rect 18656 5516 18662 5568
rect 552 5466 19412 5488
rect 552 5414 2755 5466
rect 2807 5414 2819 5466
rect 2871 5414 2883 5466
rect 2935 5414 2947 5466
rect 2999 5414 3011 5466
rect 3063 5414 7470 5466
rect 7522 5414 7534 5466
rect 7586 5414 7598 5466
rect 7650 5414 7662 5466
rect 7714 5414 7726 5466
rect 7778 5414 12185 5466
rect 12237 5414 12249 5466
rect 12301 5414 12313 5466
rect 12365 5414 12377 5466
rect 12429 5414 12441 5466
rect 12493 5414 16900 5466
rect 16952 5414 16964 5466
rect 17016 5414 17028 5466
rect 17080 5414 17092 5466
rect 17144 5414 17156 5466
rect 17208 5414 19412 5466
rect 552 5392 19412 5414
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11112 5188 11161 5216
rect 11112 5176 11118 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 11405 5151 11463 5157
rect 11405 5148 11417 5151
rect 11296 5120 11417 5148
rect 11296 5108 11302 5120
rect 11405 5117 11417 5120
rect 11451 5117 11463 5151
rect 11405 5111 11463 5117
rect 12529 5015 12587 5021
rect 12529 4981 12541 5015
rect 12575 5012 12587 5015
rect 13630 5012 13636 5024
rect 12575 4984 13636 5012
rect 12575 4981 12587 4984
rect 12529 4975 12587 4981
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 552 4922 19571 4944
rect 552 4870 5112 4922
rect 5164 4870 5176 4922
rect 5228 4870 5240 4922
rect 5292 4870 5304 4922
rect 5356 4870 5368 4922
rect 5420 4870 9827 4922
rect 9879 4870 9891 4922
rect 9943 4870 9955 4922
rect 10007 4870 10019 4922
rect 10071 4870 10083 4922
rect 10135 4870 14542 4922
rect 14594 4870 14606 4922
rect 14658 4870 14670 4922
rect 14722 4870 14734 4922
rect 14786 4870 14798 4922
rect 14850 4870 19257 4922
rect 19309 4870 19321 4922
rect 19373 4870 19385 4922
rect 19437 4870 19449 4922
rect 19501 4870 19513 4922
rect 19565 4870 19571 4922
rect 552 4848 19571 4870
rect 552 4378 19412 4400
rect 552 4326 2755 4378
rect 2807 4326 2819 4378
rect 2871 4326 2883 4378
rect 2935 4326 2947 4378
rect 2999 4326 3011 4378
rect 3063 4326 7470 4378
rect 7522 4326 7534 4378
rect 7586 4326 7598 4378
rect 7650 4326 7662 4378
rect 7714 4326 7726 4378
rect 7778 4326 12185 4378
rect 12237 4326 12249 4378
rect 12301 4326 12313 4378
rect 12365 4326 12377 4378
rect 12429 4326 12441 4378
rect 12493 4326 16900 4378
rect 16952 4326 16964 4378
rect 17016 4326 17028 4378
rect 17080 4326 17092 4378
rect 17144 4326 17156 4378
rect 17208 4326 19412 4378
rect 552 4304 19412 4326
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 8478 4128 8484 4140
rect 3752 4100 8484 4128
rect 3752 4088 3758 4100
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 552 3834 19571 3856
rect 552 3782 5112 3834
rect 5164 3782 5176 3834
rect 5228 3782 5240 3834
rect 5292 3782 5304 3834
rect 5356 3782 5368 3834
rect 5420 3782 9827 3834
rect 9879 3782 9891 3834
rect 9943 3782 9955 3834
rect 10007 3782 10019 3834
rect 10071 3782 10083 3834
rect 10135 3782 14542 3834
rect 14594 3782 14606 3834
rect 14658 3782 14670 3834
rect 14722 3782 14734 3834
rect 14786 3782 14798 3834
rect 14850 3782 19257 3834
rect 19309 3782 19321 3834
rect 19373 3782 19385 3834
rect 19437 3782 19449 3834
rect 19501 3782 19513 3834
rect 19565 3782 19571 3834
rect 552 3760 19571 3782
rect 1210 3476 1216 3528
rect 1268 3516 1274 3528
rect 6546 3516 6552 3528
rect 1268 3488 6552 3516
rect 1268 3476 1274 3488
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 552 3290 19412 3312
rect 552 3238 2755 3290
rect 2807 3238 2819 3290
rect 2871 3238 2883 3290
rect 2935 3238 2947 3290
rect 2999 3238 3011 3290
rect 3063 3238 7470 3290
rect 7522 3238 7534 3290
rect 7586 3238 7598 3290
rect 7650 3238 7662 3290
rect 7714 3238 7726 3290
rect 7778 3238 12185 3290
rect 12237 3238 12249 3290
rect 12301 3238 12313 3290
rect 12365 3238 12377 3290
rect 12429 3238 12441 3290
rect 12493 3238 16900 3290
rect 16952 3238 16964 3290
rect 17016 3238 17028 3290
rect 17080 3238 17092 3290
rect 17144 3238 17156 3290
rect 17208 3238 19412 3290
rect 552 3216 19412 3238
rect 552 2746 19571 2768
rect 552 2694 5112 2746
rect 5164 2694 5176 2746
rect 5228 2694 5240 2746
rect 5292 2694 5304 2746
rect 5356 2694 5368 2746
rect 5420 2694 9827 2746
rect 9879 2694 9891 2746
rect 9943 2694 9955 2746
rect 10007 2694 10019 2746
rect 10071 2694 10083 2746
rect 10135 2694 14542 2746
rect 14594 2694 14606 2746
rect 14658 2694 14670 2746
rect 14722 2694 14734 2746
rect 14786 2694 14798 2746
rect 14850 2694 19257 2746
rect 19309 2694 19321 2746
rect 19373 2694 19385 2746
rect 19437 2694 19449 2746
rect 19501 2694 19513 2746
rect 19565 2694 19571 2746
rect 552 2672 19571 2694
rect 552 2202 19412 2224
rect 552 2150 2755 2202
rect 2807 2150 2819 2202
rect 2871 2150 2883 2202
rect 2935 2150 2947 2202
rect 2999 2150 3011 2202
rect 3063 2150 7470 2202
rect 7522 2150 7534 2202
rect 7586 2150 7598 2202
rect 7650 2150 7662 2202
rect 7714 2150 7726 2202
rect 7778 2150 12185 2202
rect 12237 2150 12249 2202
rect 12301 2150 12313 2202
rect 12365 2150 12377 2202
rect 12429 2150 12441 2202
rect 12493 2150 16900 2202
rect 16952 2150 16964 2202
rect 17016 2150 17028 2202
rect 17080 2150 17092 2202
rect 17144 2150 17156 2202
rect 17208 2150 19412 2202
rect 552 2128 19412 2150
rect 552 1658 19571 1680
rect 552 1606 5112 1658
rect 5164 1606 5176 1658
rect 5228 1606 5240 1658
rect 5292 1606 5304 1658
rect 5356 1606 5368 1658
rect 5420 1606 9827 1658
rect 9879 1606 9891 1658
rect 9943 1606 9955 1658
rect 10007 1606 10019 1658
rect 10071 1606 10083 1658
rect 10135 1606 14542 1658
rect 14594 1606 14606 1658
rect 14658 1606 14670 1658
rect 14722 1606 14734 1658
rect 14786 1606 14798 1658
rect 14850 1606 19257 1658
rect 19309 1606 19321 1658
rect 19373 1606 19385 1658
rect 19437 1606 19449 1658
rect 19501 1606 19513 1658
rect 19565 1606 19571 1658
rect 552 1584 19571 1606
rect 552 1114 19412 1136
rect 552 1062 2755 1114
rect 2807 1062 2819 1114
rect 2871 1062 2883 1114
rect 2935 1062 2947 1114
rect 2999 1062 3011 1114
rect 3063 1062 7470 1114
rect 7522 1062 7534 1114
rect 7586 1062 7598 1114
rect 7650 1062 7662 1114
rect 7714 1062 7726 1114
rect 7778 1062 12185 1114
rect 12237 1062 12249 1114
rect 12301 1062 12313 1114
rect 12365 1062 12377 1114
rect 12429 1062 12441 1114
rect 12493 1062 16900 1114
rect 16952 1062 16964 1114
rect 17016 1062 17028 1114
rect 17080 1062 17092 1114
rect 17144 1062 17156 1114
rect 17208 1062 19412 1114
rect 552 1040 19412 1062
rect 552 570 19571 592
rect 552 518 5112 570
rect 5164 518 5176 570
rect 5228 518 5240 570
rect 5292 518 5304 570
rect 5356 518 5368 570
rect 5420 518 9827 570
rect 9879 518 9891 570
rect 9943 518 9955 570
rect 10007 518 10019 570
rect 10071 518 10083 570
rect 10135 518 14542 570
rect 14594 518 14606 570
rect 14658 518 14670 570
rect 14722 518 14734 570
rect 14786 518 14798 570
rect 14850 518 19257 570
rect 19309 518 19321 570
rect 19373 518 19385 570
rect 19437 518 19449 570
rect 19501 518 19513 570
rect 19565 518 19571 570
rect 552 496 19571 518
<< via1 >>
rect 5112 19014 5164 19066
rect 5176 19014 5228 19066
rect 5240 19014 5292 19066
rect 5304 19014 5356 19066
rect 5368 19014 5420 19066
rect 9827 19014 9879 19066
rect 9891 19014 9943 19066
rect 9955 19014 10007 19066
rect 10019 19014 10071 19066
rect 10083 19014 10135 19066
rect 14542 19014 14594 19066
rect 14606 19014 14658 19066
rect 14670 19014 14722 19066
rect 14734 19014 14786 19066
rect 14798 19014 14850 19066
rect 19257 19014 19309 19066
rect 19321 19014 19373 19066
rect 19385 19014 19437 19066
rect 19449 19014 19501 19066
rect 19513 19014 19565 19066
rect 8668 18912 8720 18964
rect 9128 18844 9180 18896
rect 848 18776 900 18828
rect 2504 18776 2556 18828
rect 4160 18776 4212 18828
rect 5816 18776 5868 18828
rect 7472 18776 7524 18828
rect 6460 18708 6512 18760
rect 10784 18776 10836 18828
rect 12440 18776 12492 18828
rect 14096 18776 14148 18828
rect 15752 18776 15804 18828
rect 17408 18776 17460 18828
rect 9220 18640 9272 18692
rect 9588 18708 9640 18760
rect 9680 18640 9732 18692
rect 7012 18572 7064 18624
rect 8576 18572 8628 18624
rect 9496 18615 9548 18624
rect 9496 18581 9505 18615
rect 9505 18581 9539 18615
rect 9539 18581 9548 18615
rect 9496 18572 9548 18581
rect 10600 18572 10652 18624
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16764 18572 16816 18624
rect 2755 18470 2807 18522
rect 2819 18470 2871 18522
rect 2883 18470 2935 18522
rect 2947 18470 2999 18522
rect 3011 18470 3063 18522
rect 7470 18470 7522 18522
rect 7534 18470 7586 18522
rect 7598 18470 7650 18522
rect 7662 18470 7714 18522
rect 7726 18470 7778 18522
rect 12185 18470 12237 18522
rect 12249 18470 12301 18522
rect 12313 18470 12365 18522
rect 12377 18470 12429 18522
rect 12441 18470 12493 18522
rect 16900 18470 16952 18522
rect 16964 18470 17016 18522
rect 17028 18470 17080 18522
rect 17092 18470 17144 18522
rect 17156 18470 17208 18522
rect 9036 18300 9088 18352
rect 7012 18232 7064 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 8300 18232 8352 18284
rect 8944 18232 8996 18284
rect 9312 18368 9364 18420
rect 3608 18207 3660 18216
rect 3608 18173 3617 18207
rect 3617 18173 3651 18207
rect 3651 18173 3660 18207
rect 3608 18164 3660 18173
rect 3792 18164 3844 18216
rect 8300 18096 8352 18148
rect 3332 18028 3384 18080
rect 4988 18028 5040 18080
rect 6736 18071 6788 18080
rect 6736 18037 6745 18071
rect 6745 18037 6779 18071
rect 6779 18037 6788 18071
rect 6736 18028 6788 18037
rect 6828 18071 6880 18080
rect 6828 18037 6837 18071
rect 6837 18037 6871 18071
rect 6871 18037 6880 18071
rect 6828 18028 6880 18037
rect 8392 18071 8444 18080
rect 8392 18037 8401 18071
rect 8401 18037 8435 18071
rect 8435 18037 8444 18071
rect 8392 18028 8444 18037
rect 9404 18164 9456 18216
rect 8944 18096 8996 18148
rect 9128 18028 9180 18080
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 16764 18207 16816 18216
rect 16764 18173 16773 18207
rect 16773 18173 16807 18207
rect 16807 18173 16816 18207
rect 16764 18164 16816 18173
rect 14464 18028 14516 18080
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 5112 17926 5164 17978
rect 5176 17926 5228 17978
rect 5240 17926 5292 17978
rect 5304 17926 5356 17978
rect 5368 17926 5420 17978
rect 9827 17926 9879 17978
rect 9891 17926 9943 17978
rect 9955 17926 10007 17978
rect 10019 17926 10071 17978
rect 10083 17926 10135 17978
rect 14542 17926 14594 17978
rect 14606 17926 14658 17978
rect 14670 17926 14722 17978
rect 14734 17926 14786 17978
rect 14798 17926 14850 17978
rect 19257 17926 19309 17978
rect 19321 17926 19373 17978
rect 19385 17926 19437 17978
rect 19449 17926 19501 17978
rect 19513 17926 19565 17978
rect 2044 17824 2096 17876
rect 4896 17824 4948 17876
rect 6736 17824 6788 17876
rect 8392 17824 8444 17876
rect 9036 17867 9088 17876
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 848 17620 900 17672
rect 2320 17688 2372 17740
rect 3792 17756 3844 17808
rect 3332 17731 3384 17740
rect 3332 17697 3366 17731
rect 3366 17697 3384 17731
rect 3332 17688 3384 17697
rect 4712 17688 4764 17740
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 6828 17688 6880 17740
rect 8392 17688 8444 17740
rect 4988 17620 5040 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 8300 17620 8352 17672
rect 9496 17731 9548 17740
rect 9496 17697 9505 17731
rect 9505 17697 9539 17731
rect 9539 17697 9548 17731
rect 9496 17688 9548 17697
rect 9680 17731 9732 17740
rect 9680 17697 9689 17731
rect 9689 17697 9723 17731
rect 9723 17697 9732 17731
rect 9680 17688 9732 17697
rect 10232 17688 10284 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 11704 17688 11756 17740
rect 14464 17799 14516 17808
rect 14464 17765 14473 17799
rect 14473 17765 14507 17799
rect 14507 17765 14516 17799
rect 14464 17756 14516 17765
rect 16672 17756 16724 17808
rect 11428 17620 11480 17672
rect 13544 17620 13596 17672
rect 7932 17552 7984 17604
rect 16120 17620 16172 17672
rect 3240 17484 3292 17536
rect 5264 17484 5316 17536
rect 5632 17484 5684 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 8392 17484 8444 17536
rect 8484 17484 8536 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 9496 17484 9548 17536
rect 10416 17484 10468 17536
rect 11428 17527 11480 17536
rect 11428 17493 11437 17527
rect 11437 17493 11471 17527
rect 11471 17493 11480 17527
rect 11428 17484 11480 17493
rect 2755 17382 2807 17434
rect 2819 17382 2871 17434
rect 2883 17382 2935 17434
rect 2947 17382 2999 17434
rect 3011 17382 3063 17434
rect 7470 17382 7522 17434
rect 7534 17382 7586 17434
rect 7598 17382 7650 17434
rect 7662 17382 7714 17434
rect 7726 17382 7778 17434
rect 12185 17382 12237 17434
rect 12249 17382 12301 17434
rect 12313 17382 12365 17434
rect 12377 17382 12429 17434
rect 12441 17382 12493 17434
rect 16900 17382 16952 17434
rect 16964 17382 17016 17434
rect 17028 17382 17080 17434
rect 17092 17382 17144 17434
rect 17156 17382 17208 17434
rect 3608 17280 3660 17332
rect 5080 17280 5132 17332
rect 5540 17280 5592 17332
rect 6736 17280 6788 17332
rect 8852 17280 8904 17332
rect 3976 17144 4028 17196
rect 6828 17212 6880 17264
rect 2044 17119 2096 17128
rect 2044 17085 2053 17119
rect 2053 17085 2087 17119
rect 2087 17085 2096 17119
rect 2044 17076 2096 17085
rect 2136 17076 2188 17128
rect 3240 17076 3292 17128
rect 4160 17076 4212 17128
rect 5080 17144 5132 17196
rect 4988 17119 5040 17128
rect 4988 17085 4998 17119
rect 4998 17085 5032 17119
rect 5032 17085 5040 17119
rect 4988 17076 5040 17085
rect 5264 17119 5316 17128
rect 5264 17085 5273 17119
rect 5273 17085 5307 17119
rect 5307 17085 5316 17119
rect 5264 17076 5316 17085
rect 5540 17076 5592 17128
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 5816 17119 5868 17128
rect 5816 17085 5823 17119
rect 5823 17085 5868 17119
rect 5816 17076 5868 17085
rect 3332 17008 3384 17060
rect 2504 16983 2556 16992
rect 2504 16949 2513 16983
rect 2513 16949 2547 16983
rect 2547 16949 2556 16983
rect 2504 16940 2556 16949
rect 5908 17051 5960 17060
rect 5908 17017 5917 17051
rect 5917 17017 5951 17051
rect 5951 17017 5960 17051
rect 5908 17008 5960 17017
rect 8208 17076 8260 17128
rect 5448 16940 5500 16992
rect 5540 16983 5592 16992
rect 5540 16949 5549 16983
rect 5549 16949 5583 16983
rect 5583 16949 5592 16983
rect 5540 16940 5592 16949
rect 5632 16940 5684 16992
rect 7196 17008 7248 17060
rect 7840 17051 7892 17060
rect 7840 17017 7858 17051
rect 7858 17017 7892 17051
rect 7840 17008 7892 17017
rect 9680 17008 9732 17060
rect 5112 16838 5164 16890
rect 5176 16838 5228 16890
rect 5240 16838 5292 16890
rect 5304 16838 5356 16890
rect 5368 16838 5420 16890
rect 9827 16838 9879 16890
rect 9891 16838 9943 16890
rect 9955 16838 10007 16890
rect 10019 16838 10071 16890
rect 10083 16838 10135 16890
rect 14542 16838 14594 16890
rect 14606 16838 14658 16890
rect 14670 16838 14722 16890
rect 14734 16838 14786 16890
rect 14798 16838 14850 16890
rect 19257 16838 19309 16890
rect 19321 16838 19373 16890
rect 19385 16838 19437 16890
rect 19449 16838 19501 16890
rect 19513 16838 19565 16890
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 3976 16779 4028 16788
rect 3976 16745 3985 16779
rect 3985 16745 4019 16779
rect 4019 16745 4028 16779
rect 3976 16736 4028 16745
rect 4988 16736 5040 16788
rect 2504 16643 2556 16652
rect 2504 16609 2513 16643
rect 2513 16609 2547 16643
rect 2547 16609 2556 16643
rect 2504 16600 2556 16609
rect 3240 16600 3292 16652
rect 5540 16600 5592 16652
rect 5632 16600 5684 16652
rect 6184 16668 6236 16720
rect 6092 16643 6144 16652
rect 6092 16609 6101 16643
rect 6101 16609 6135 16643
rect 6135 16609 6144 16643
rect 6092 16600 6144 16609
rect 6460 16736 6512 16788
rect 6828 16736 6880 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 5264 16575 5316 16584
rect 5264 16541 5273 16575
rect 5273 16541 5307 16575
rect 5307 16541 5316 16575
rect 5264 16532 5316 16541
rect 6644 16600 6696 16652
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 8760 16668 8812 16720
rect 9680 16736 9732 16788
rect 7932 16600 7984 16652
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 8392 16600 8444 16652
rect 9956 16711 10008 16720
rect 9956 16677 9965 16711
rect 9965 16677 9999 16711
rect 9999 16677 10008 16711
rect 9956 16668 10008 16677
rect 11520 16736 11572 16788
rect 11428 16668 11480 16720
rect 9220 16600 9272 16652
rect 7104 16464 7156 16516
rect 9128 16464 9180 16516
rect 9680 16532 9732 16584
rect 10232 16600 10284 16652
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 11244 16600 11296 16652
rect 11796 16643 11848 16652
rect 11796 16609 11805 16643
rect 11805 16609 11839 16643
rect 11839 16609 11848 16643
rect 11796 16600 11848 16609
rect 12072 16600 12124 16652
rect 9588 16464 9640 16516
rect 11980 16532 12032 16584
rect 5448 16396 5500 16448
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 8852 16439 8904 16448
rect 8852 16405 8861 16439
rect 8861 16405 8895 16439
rect 8895 16405 8904 16439
rect 8852 16396 8904 16405
rect 8944 16396 8996 16448
rect 10876 16396 10928 16448
rect 11612 16396 11664 16448
rect 11796 16396 11848 16448
rect 11980 16396 12032 16448
rect 12624 16532 12676 16584
rect 15200 16532 15252 16584
rect 2755 16294 2807 16346
rect 2819 16294 2871 16346
rect 2883 16294 2935 16346
rect 2947 16294 2999 16346
rect 3011 16294 3063 16346
rect 7470 16294 7522 16346
rect 7534 16294 7586 16346
rect 7598 16294 7650 16346
rect 7662 16294 7714 16346
rect 7726 16294 7778 16346
rect 12185 16294 12237 16346
rect 12249 16294 12301 16346
rect 12313 16294 12365 16346
rect 12377 16294 12429 16346
rect 12441 16294 12493 16346
rect 16900 16294 16952 16346
rect 16964 16294 17016 16346
rect 17028 16294 17080 16346
rect 17092 16294 17144 16346
rect 17156 16294 17208 16346
rect 5264 16192 5316 16244
rect 6276 16192 6328 16244
rect 8484 16192 8536 16244
rect 9220 16192 9272 16244
rect 2136 16124 2188 16176
rect 10508 16192 10560 16244
rect 1768 16056 1820 16108
rect 9404 16167 9456 16176
rect 9404 16133 9413 16167
rect 9413 16133 9447 16167
rect 9447 16133 9456 16167
rect 9404 16124 9456 16133
rect 7104 16099 7156 16108
rect 7104 16065 7113 16099
rect 7113 16065 7147 16099
rect 7147 16065 7156 16099
rect 7104 16056 7156 16065
rect 8760 16099 8812 16108
rect 8760 16065 8769 16099
rect 8769 16065 8803 16099
rect 8803 16065 8812 16099
rect 8760 16056 8812 16065
rect 10876 16192 10928 16244
rect 12532 16192 12584 16244
rect 2136 16031 2188 16040
rect 2136 15997 2145 16031
rect 2145 15997 2179 16031
rect 2179 15997 2188 16031
rect 2136 15988 2188 15997
rect 2412 15988 2464 16040
rect 8024 15988 8076 16040
rect 8944 15988 8996 16040
rect 9036 16031 9088 16040
rect 9036 15997 9045 16031
rect 9045 15997 9079 16031
rect 9079 15997 9088 16031
rect 9036 15988 9088 15997
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 9588 16031 9640 16040
rect 9588 15997 9597 16031
rect 9597 15997 9631 16031
rect 9631 15997 9640 16031
rect 9588 15988 9640 15997
rect 2228 15920 2280 15972
rect 2504 15963 2556 15972
rect 2504 15929 2513 15963
rect 2513 15929 2547 15963
rect 2547 15929 2556 15963
rect 2504 15920 2556 15929
rect 10600 15988 10652 16040
rect 11244 15988 11296 16040
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 11612 16031 11664 16040
rect 11612 15997 11621 16031
rect 11621 15997 11655 16031
rect 11655 15997 11664 16031
rect 11612 15988 11664 15997
rect 12532 15988 12584 16040
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 10416 15920 10468 15972
rect 1308 15852 1360 15904
rect 3240 15852 3292 15904
rect 6828 15895 6880 15904
rect 6828 15861 6837 15895
rect 6837 15861 6871 15895
rect 6871 15861 6880 15895
rect 6828 15852 6880 15861
rect 7840 15852 7892 15904
rect 8484 15895 8536 15904
rect 8484 15861 8493 15895
rect 8493 15861 8527 15895
rect 8527 15861 8536 15895
rect 8484 15852 8536 15861
rect 12256 15852 12308 15904
rect 14832 15852 14884 15904
rect 15200 15852 15252 15904
rect 5112 15750 5164 15802
rect 5176 15750 5228 15802
rect 5240 15750 5292 15802
rect 5304 15750 5356 15802
rect 5368 15750 5420 15802
rect 9827 15750 9879 15802
rect 9891 15750 9943 15802
rect 9955 15750 10007 15802
rect 10019 15750 10071 15802
rect 10083 15750 10135 15802
rect 14542 15750 14594 15802
rect 14606 15750 14658 15802
rect 14670 15750 14722 15802
rect 14734 15750 14786 15802
rect 14798 15750 14850 15802
rect 19257 15750 19309 15802
rect 19321 15750 19373 15802
rect 19385 15750 19437 15802
rect 19449 15750 19501 15802
rect 19513 15750 19565 15802
rect 2136 15648 2188 15700
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 1768 15623 1820 15632
rect 1768 15589 1777 15623
rect 1777 15589 1811 15623
rect 1811 15589 1820 15623
rect 1768 15580 1820 15589
rect 2228 15580 2280 15632
rect 3332 15648 3384 15700
rect 10508 15691 10560 15700
rect 10508 15657 10517 15691
rect 10517 15657 10551 15691
rect 10551 15657 10560 15691
rect 10508 15648 10560 15657
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 13820 15648 13872 15700
rect 9404 15623 9456 15632
rect 9404 15589 9438 15623
rect 9438 15589 9456 15623
rect 9404 15580 9456 15589
rect 1952 15444 2004 15496
rect 2504 15444 2556 15496
rect 3516 15555 3568 15564
rect 3516 15521 3534 15555
rect 3534 15521 3568 15555
rect 3516 15512 3568 15521
rect 3792 15555 3844 15564
rect 3792 15521 3801 15555
rect 3801 15521 3835 15555
rect 3835 15521 3844 15555
rect 3792 15512 3844 15521
rect 7196 15512 7248 15564
rect 8668 15555 8720 15564
rect 8668 15521 8677 15555
rect 8677 15521 8711 15555
rect 8711 15521 8720 15555
rect 8668 15512 8720 15521
rect 9220 15512 9272 15564
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 11152 15555 11204 15564
rect 11152 15521 11161 15555
rect 11161 15521 11195 15555
rect 11195 15521 11204 15555
rect 11152 15512 11204 15521
rect 11704 15512 11756 15564
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 11980 15555 12032 15564
rect 11980 15521 11989 15555
rect 11989 15521 12023 15555
rect 12023 15521 12032 15555
rect 11980 15512 12032 15521
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 2596 15376 2648 15428
rect 11152 15376 11204 15428
rect 1032 15351 1084 15360
rect 1032 15317 1041 15351
rect 1041 15317 1075 15351
rect 1075 15317 1084 15351
rect 1032 15308 1084 15317
rect 1308 15351 1360 15360
rect 1308 15317 1317 15351
rect 1317 15317 1351 15351
rect 1351 15317 1360 15351
rect 1308 15308 1360 15317
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 10600 15308 10652 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 2755 15206 2807 15258
rect 2819 15206 2871 15258
rect 2883 15206 2935 15258
rect 2947 15206 2999 15258
rect 3011 15206 3063 15258
rect 7470 15206 7522 15258
rect 7534 15206 7586 15258
rect 7598 15206 7650 15258
rect 7662 15206 7714 15258
rect 7726 15206 7778 15258
rect 12185 15206 12237 15258
rect 12249 15206 12301 15258
rect 12313 15206 12365 15258
rect 12377 15206 12429 15258
rect 12441 15206 12493 15258
rect 16900 15206 16952 15258
rect 16964 15206 17016 15258
rect 17028 15206 17080 15258
rect 17092 15206 17144 15258
rect 17156 15206 17208 15258
rect 3240 15104 3292 15156
rect 3516 15104 3568 15156
rect 9036 15104 9088 15156
rect 11520 15147 11572 15156
rect 11520 15113 11529 15147
rect 11529 15113 11563 15147
rect 11563 15113 11572 15147
rect 11520 15104 11572 15113
rect 12900 15104 12952 15156
rect 848 15011 900 15020
rect 848 14977 857 15011
rect 857 14977 891 15011
rect 891 14977 900 15011
rect 848 14968 900 14977
rect 1032 14832 1084 14884
rect 2320 14900 2372 14952
rect 4160 14900 4212 14952
rect 4804 14900 4856 14952
rect 5816 14900 5868 14952
rect 6276 14943 6328 14952
rect 6276 14909 6285 14943
rect 6285 14909 6319 14943
rect 6319 14909 6328 14943
rect 6276 14900 6328 14909
rect 6828 14900 6880 14952
rect 9128 14900 9180 14952
rect 4528 14832 4580 14884
rect 8944 14832 8996 14884
rect 10600 14832 10652 14884
rect 11612 14832 11664 14884
rect 11888 14832 11940 14884
rect 14924 14943 14976 14952
rect 14924 14909 14933 14943
rect 14933 14909 14967 14943
rect 14967 14909 14976 14943
rect 14924 14900 14976 14909
rect 15200 14832 15252 14884
rect 16212 14832 16264 14884
rect 2228 14807 2280 14816
rect 2228 14773 2237 14807
rect 2237 14773 2271 14807
rect 2271 14773 2280 14807
rect 2228 14764 2280 14773
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 4160 14764 4212 14816
rect 4988 14764 5040 14816
rect 7288 14764 7340 14816
rect 15476 14807 15528 14816
rect 15476 14773 15485 14807
rect 15485 14773 15519 14807
rect 15519 14773 15528 14807
rect 15476 14764 15528 14773
rect 5112 14662 5164 14714
rect 5176 14662 5228 14714
rect 5240 14662 5292 14714
rect 5304 14662 5356 14714
rect 5368 14662 5420 14714
rect 9827 14662 9879 14714
rect 9891 14662 9943 14714
rect 9955 14662 10007 14714
rect 10019 14662 10071 14714
rect 10083 14662 10135 14714
rect 14542 14662 14594 14714
rect 14606 14662 14658 14714
rect 14670 14662 14722 14714
rect 14734 14662 14786 14714
rect 14798 14662 14850 14714
rect 19257 14662 19309 14714
rect 19321 14662 19373 14714
rect 19385 14662 19437 14714
rect 19449 14662 19501 14714
rect 19513 14662 19565 14714
rect 1768 14560 1820 14612
rect 2228 14492 2280 14544
rect 2872 14492 2924 14544
rect 4068 14492 4120 14544
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 8484 14560 8536 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 5080 14492 5132 14544
rect 11428 14492 11480 14544
rect 12072 14492 12124 14544
rect 5540 14424 5592 14476
rect 7104 14424 7156 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 7288 14467 7340 14476
rect 7288 14433 7297 14467
rect 7297 14433 7331 14467
rect 7331 14433 7340 14467
rect 7288 14424 7340 14433
rect 5448 14356 5500 14408
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 15292 14492 15344 14544
rect 1952 14331 2004 14340
rect 1952 14297 1961 14331
rect 1961 14297 1995 14331
rect 1995 14297 2004 14331
rect 1952 14288 2004 14297
rect 5172 14288 5224 14340
rect 11888 14399 11940 14408
rect 11888 14365 11897 14399
rect 11897 14365 11931 14399
rect 11931 14365 11940 14399
rect 11888 14356 11940 14365
rect 8760 14288 8812 14340
rect 10784 14288 10836 14340
rect 11704 14331 11756 14340
rect 11704 14297 11713 14331
rect 11713 14297 11747 14331
rect 11747 14297 11756 14331
rect 12532 14424 12584 14476
rect 12716 14467 12768 14476
rect 12716 14433 12750 14467
rect 12750 14433 12768 14467
rect 12716 14424 12768 14433
rect 14924 14467 14976 14476
rect 14924 14433 14933 14467
rect 14933 14433 14967 14467
rect 14967 14433 14976 14467
rect 14924 14424 14976 14433
rect 15108 14424 15160 14476
rect 11704 14288 11756 14297
rect 2136 14263 2188 14272
rect 2136 14229 2145 14263
rect 2145 14229 2179 14263
rect 2179 14229 2188 14263
rect 2136 14220 2188 14229
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4620 14263 4672 14272
rect 4620 14229 4629 14263
rect 4629 14229 4663 14263
rect 4663 14229 4672 14263
rect 4620 14220 4672 14229
rect 4988 14220 5040 14272
rect 5356 14220 5408 14272
rect 8392 14220 8444 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 12808 14220 12860 14272
rect 13820 14263 13872 14272
rect 13820 14229 13829 14263
rect 13829 14229 13863 14263
rect 13863 14229 13872 14263
rect 13820 14220 13872 14229
rect 2755 14118 2807 14170
rect 2819 14118 2871 14170
rect 2883 14118 2935 14170
rect 2947 14118 2999 14170
rect 3011 14118 3063 14170
rect 7470 14118 7522 14170
rect 7534 14118 7586 14170
rect 7598 14118 7650 14170
rect 7662 14118 7714 14170
rect 7726 14118 7778 14170
rect 12185 14118 12237 14170
rect 12249 14118 12301 14170
rect 12313 14118 12365 14170
rect 12377 14118 12429 14170
rect 12441 14118 12493 14170
rect 16900 14118 16952 14170
rect 16964 14118 17016 14170
rect 17028 14118 17080 14170
rect 17092 14118 17144 14170
rect 17156 14118 17208 14170
rect 4344 14016 4396 14068
rect 1308 13812 1360 13864
rect 2780 13880 2832 13932
rect 4804 13948 4856 14000
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 4620 13812 4672 13864
rect 5540 14059 5592 14068
rect 5540 14025 5549 14059
rect 5549 14025 5583 14059
rect 5583 14025 5592 14059
rect 5540 14016 5592 14025
rect 11704 14016 11756 14068
rect 12072 14059 12124 14068
rect 12072 14025 12081 14059
rect 12081 14025 12115 14059
rect 12115 14025 12124 14059
rect 12072 14016 12124 14025
rect 12716 14016 12768 14068
rect 5816 13948 5868 14000
rect 5632 13880 5684 13932
rect 6276 13880 6328 13932
rect 7288 13948 7340 14000
rect 6920 13923 6972 13932
rect 6920 13889 6929 13923
rect 6929 13889 6963 13923
rect 6963 13889 6972 13923
rect 6920 13880 6972 13889
rect 4344 13744 4396 13796
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 5448 13812 5500 13864
rect 8392 13812 8444 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 11060 13787 11112 13796
rect 11060 13753 11069 13787
rect 11069 13753 11103 13787
rect 11103 13753 11112 13787
rect 11060 13744 11112 13753
rect 11520 13744 11572 13796
rect 12624 13812 12676 13864
rect 12808 13812 12860 13864
rect 13820 13812 13872 13864
rect 15108 13812 15160 13864
rect 16212 13855 16264 13864
rect 16212 13821 16221 13855
rect 16221 13821 16255 13855
rect 16255 13821 16264 13855
rect 16212 13812 16264 13821
rect 16488 13855 16540 13864
rect 16488 13821 16497 13855
rect 16497 13821 16531 13855
rect 16531 13821 16540 13855
rect 16488 13812 16540 13821
rect 15936 13744 15988 13796
rect 5172 13719 5224 13728
rect 5172 13685 5181 13719
rect 5181 13685 5215 13719
rect 5215 13685 5224 13719
rect 5172 13676 5224 13685
rect 5448 13676 5500 13728
rect 10232 13676 10284 13728
rect 10876 13676 10928 13728
rect 11796 13676 11848 13728
rect 5112 13574 5164 13626
rect 5176 13574 5228 13626
rect 5240 13574 5292 13626
rect 5304 13574 5356 13626
rect 5368 13574 5420 13626
rect 9827 13574 9879 13626
rect 9891 13574 9943 13626
rect 9955 13574 10007 13626
rect 10019 13574 10071 13626
rect 10083 13574 10135 13626
rect 14542 13574 14594 13626
rect 14606 13574 14658 13626
rect 14670 13574 14722 13626
rect 14734 13574 14786 13626
rect 14798 13574 14850 13626
rect 19257 13574 19309 13626
rect 19321 13574 19373 13626
rect 19385 13574 19437 13626
rect 19449 13574 19501 13626
rect 19513 13574 19565 13626
rect 2320 13472 2372 13524
rect 5080 13472 5132 13524
rect 11152 13472 11204 13524
rect 1308 13447 1360 13456
rect 1308 13413 1342 13447
rect 1342 13413 1360 13447
rect 1308 13404 1360 13413
rect 4068 13404 4120 13456
rect 7840 13404 7892 13456
rect 9036 13404 9088 13456
rect 9404 13404 9456 13456
rect 2044 13336 2096 13388
rect 2504 13379 2556 13388
rect 2504 13345 2513 13379
rect 2513 13345 2547 13379
rect 2547 13345 2556 13379
rect 2504 13336 2556 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3148 13336 3200 13388
rect 5448 13336 5500 13388
rect 6920 13336 6972 13388
rect 9128 13336 9180 13388
rect 9956 13336 10008 13388
rect 4712 13268 4764 13320
rect 4436 13200 4488 13252
rect 8300 13311 8352 13320
rect 8300 13277 8309 13311
rect 8309 13277 8343 13311
rect 8343 13277 8352 13311
rect 8300 13268 8352 13277
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 11980 13379 12032 13388
rect 11980 13345 11989 13379
rect 11989 13345 12023 13379
rect 12023 13345 12032 13379
rect 11980 13336 12032 13345
rect 15016 13472 15068 13524
rect 16488 13472 16540 13524
rect 15108 13379 15160 13388
rect 15108 13345 15117 13379
rect 15117 13345 15151 13379
rect 15151 13345 15160 13379
rect 15108 13336 15160 13345
rect 16212 13379 16264 13388
rect 16212 13345 16221 13379
rect 16221 13345 16255 13379
rect 16255 13345 16264 13379
rect 16212 13336 16264 13345
rect 16488 13336 16540 13388
rect 11336 13200 11388 13252
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 1768 13132 1820 13184
rect 2964 13132 3016 13184
rect 3976 13132 4028 13184
rect 6092 13132 6144 13184
rect 10968 13175 11020 13184
rect 10968 13141 10977 13175
rect 10977 13141 11011 13175
rect 11011 13141 11020 13175
rect 10968 13132 11020 13141
rect 13728 13132 13780 13184
rect 15200 13132 15252 13184
rect 17868 13175 17920 13184
rect 17868 13141 17877 13175
rect 17877 13141 17911 13175
rect 17911 13141 17920 13175
rect 17868 13132 17920 13141
rect 2755 13030 2807 13082
rect 2819 13030 2871 13082
rect 2883 13030 2935 13082
rect 2947 13030 2999 13082
rect 3011 13030 3063 13082
rect 7470 13030 7522 13082
rect 7534 13030 7586 13082
rect 7598 13030 7650 13082
rect 7662 13030 7714 13082
rect 7726 13030 7778 13082
rect 12185 13030 12237 13082
rect 12249 13030 12301 13082
rect 12313 13030 12365 13082
rect 12377 13030 12429 13082
rect 12441 13030 12493 13082
rect 16900 13030 16952 13082
rect 16964 13030 17016 13082
rect 17028 13030 17080 13082
rect 17092 13030 17144 13082
rect 17156 13030 17208 13082
rect 2780 12928 2832 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 8300 12928 8352 12980
rect 8116 12860 8168 12912
rect 9680 12928 9732 12980
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 8668 12860 8720 12912
rect 10692 12860 10744 12912
rect 11060 12928 11112 12980
rect 12072 12928 12124 12980
rect 12532 12928 12584 12980
rect 11704 12860 11756 12912
rect 2504 12792 2556 12844
rect 1768 12724 1820 12776
rect 2596 12724 2648 12776
rect 4712 12792 4764 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 2688 12588 2740 12640
rect 3976 12699 4028 12708
rect 3976 12665 3985 12699
rect 3985 12665 4019 12699
rect 4019 12665 4028 12699
rect 3976 12656 4028 12665
rect 3148 12588 3200 12640
rect 5448 12724 5500 12776
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7840 12724 7892 12776
rect 9036 12792 9088 12844
rect 10968 12792 11020 12844
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 8944 12724 8996 12776
rect 9404 12724 9456 12776
rect 9680 12724 9732 12776
rect 10232 12724 10284 12776
rect 10324 12724 10376 12776
rect 4620 12656 4672 12708
rect 4896 12588 4948 12640
rect 5448 12588 5500 12640
rect 7104 12588 7156 12640
rect 8944 12588 8996 12640
rect 9404 12588 9456 12640
rect 10232 12588 10284 12640
rect 10876 12724 10928 12776
rect 11336 12767 11388 12776
rect 11336 12733 11345 12767
rect 11345 12733 11379 12767
rect 11379 12733 11388 12767
rect 11336 12724 11388 12733
rect 15016 12724 15068 12776
rect 15108 12767 15160 12776
rect 15108 12733 15117 12767
rect 15117 12733 15151 12767
rect 15151 12733 15160 12767
rect 15108 12724 15160 12733
rect 10968 12656 11020 12708
rect 11520 12699 11572 12708
rect 11520 12665 11529 12699
rect 11529 12665 11563 12699
rect 11563 12665 11572 12699
rect 11520 12656 11572 12665
rect 13360 12656 13412 12708
rect 16304 12656 16356 12708
rect 5112 12486 5164 12538
rect 5176 12486 5228 12538
rect 5240 12486 5292 12538
rect 5304 12486 5356 12538
rect 5368 12486 5420 12538
rect 9827 12486 9879 12538
rect 9891 12486 9943 12538
rect 9955 12486 10007 12538
rect 10019 12486 10071 12538
rect 10083 12486 10135 12538
rect 14542 12486 14594 12538
rect 14606 12486 14658 12538
rect 14670 12486 14722 12538
rect 14734 12486 14786 12538
rect 14798 12486 14850 12538
rect 19257 12486 19309 12538
rect 19321 12486 19373 12538
rect 19385 12486 19437 12538
rect 19449 12486 19501 12538
rect 19513 12486 19565 12538
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 4988 12384 5040 12436
rect 2780 12359 2832 12368
rect 2780 12325 2789 12359
rect 2789 12325 2823 12359
rect 2823 12325 2832 12359
rect 2780 12316 2832 12325
rect 3240 12316 3292 12368
rect 2504 12248 2556 12300
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 4252 12248 4304 12300
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 5632 12316 5684 12368
rect 4804 12248 4856 12257
rect 7104 12248 7156 12300
rect 10140 12316 10192 12368
rect 10968 12384 11020 12436
rect 12624 12384 12676 12436
rect 9404 12248 9456 12300
rect 12072 12316 12124 12368
rect 14464 12316 14516 12368
rect 15016 12316 15068 12368
rect 11060 12248 11112 12300
rect 3056 12180 3108 12232
rect 3332 12180 3384 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 6092 12180 6144 12232
rect 8484 12180 8536 12232
rect 9772 12180 9824 12232
rect 10232 12180 10284 12232
rect 2688 12044 2740 12096
rect 3148 12044 3200 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4068 12044 4120 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 9864 12112 9916 12164
rect 10876 12180 10928 12232
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 13728 12248 13780 12300
rect 7196 12044 7248 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 10876 12044 10928 12096
rect 2755 11942 2807 11994
rect 2819 11942 2871 11994
rect 2883 11942 2935 11994
rect 2947 11942 2999 11994
rect 3011 11942 3063 11994
rect 7470 11942 7522 11994
rect 7534 11942 7586 11994
rect 7598 11942 7650 11994
rect 7662 11942 7714 11994
rect 7726 11942 7778 11994
rect 12185 11942 12237 11994
rect 12249 11942 12301 11994
rect 12313 11942 12365 11994
rect 12377 11942 12429 11994
rect 12441 11942 12493 11994
rect 16900 11942 16952 11994
rect 16964 11942 17016 11994
rect 17028 11942 17080 11994
rect 17092 11942 17144 11994
rect 17156 11942 17208 11994
rect 3148 11840 3200 11892
rect 4896 11883 4948 11892
rect 4896 11849 4905 11883
rect 4905 11849 4939 11883
rect 4939 11849 4948 11883
rect 4896 11840 4948 11849
rect 4712 11772 4764 11824
rect 7840 11840 7892 11892
rect 11060 11840 11112 11892
rect 15200 11840 15252 11892
rect 15384 11840 15436 11892
rect 15936 11840 15988 11892
rect 2964 11704 3016 11756
rect 3240 11704 3292 11756
rect 2504 11679 2556 11688
rect 2504 11645 2513 11679
rect 2513 11645 2547 11679
rect 2547 11645 2556 11679
rect 2504 11636 2556 11645
rect 2596 11636 2648 11688
rect 5632 11704 5684 11756
rect 5816 11704 5868 11756
rect 13452 11772 13504 11824
rect 16672 11772 16724 11824
rect 3056 11568 3108 11620
rect 3976 11568 4028 11620
rect 6092 11679 6144 11688
rect 6092 11645 6101 11679
rect 6101 11645 6135 11679
rect 6135 11645 6144 11679
rect 6092 11636 6144 11645
rect 3332 11500 3384 11552
rect 5448 11500 5500 11552
rect 6000 11500 6052 11552
rect 8392 11704 8444 11756
rect 10140 11704 10192 11756
rect 14464 11704 14516 11756
rect 15752 11704 15804 11756
rect 16764 11704 16816 11756
rect 8300 11636 8352 11688
rect 9772 11636 9824 11688
rect 10600 11679 10652 11688
rect 10600 11645 10609 11679
rect 10609 11645 10643 11679
rect 10643 11645 10652 11679
rect 10600 11636 10652 11645
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 12624 11636 12676 11688
rect 13360 11636 13412 11688
rect 13728 11636 13780 11688
rect 15200 11679 15252 11688
rect 15200 11645 15209 11679
rect 15209 11645 15243 11679
rect 15243 11645 15252 11679
rect 15200 11636 15252 11645
rect 15292 11636 15344 11688
rect 16028 11636 16080 11688
rect 16304 11636 16356 11688
rect 6644 11568 6696 11620
rect 8852 11568 8904 11620
rect 9864 11568 9916 11620
rect 14188 11568 14240 11620
rect 14924 11568 14976 11620
rect 9588 11500 9640 11552
rect 10416 11500 10468 11552
rect 10600 11500 10652 11552
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 15476 11500 15528 11552
rect 16396 11500 16448 11552
rect 16856 11500 16908 11552
rect 5112 11398 5164 11450
rect 5176 11398 5228 11450
rect 5240 11398 5292 11450
rect 5304 11398 5356 11450
rect 5368 11398 5420 11450
rect 9827 11398 9879 11450
rect 9891 11398 9943 11450
rect 9955 11398 10007 11450
rect 10019 11398 10071 11450
rect 10083 11398 10135 11450
rect 14542 11398 14594 11450
rect 14606 11398 14658 11450
rect 14670 11398 14722 11450
rect 14734 11398 14786 11450
rect 14798 11398 14850 11450
rect 19257 11398 19309 11450
rect 19321 11398 19373 11450
rect 19385 11398 19437 11450
rect 19449 11398 19501 11450
rect 19513 11398 19565 11450
rect 3148 11296 3200 11348
rect 4068 11339 4120 11348
rect 4068 11305 4077 11339
rect 4077 11305 4111 11339
rect 4111 11305 4120 11339
rect 4068 11296 4120 11305
rect 4252 11339 4304 11348
rect 4252 11305 4261 11339
rect 4261 11305 4295 11339
rect 4295 11305 4304 11339
rect 4252 11296 4304 11305
rect 6092 11296 6144 11348
rect 6644 11339 6696 11348
rect 6644 11305 6653 11339
rect 6653 11305 6687 11339
rect 6687 11305 6696 11339
rect 6644 11296 6696 11305
rect 8392 11296 8444 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 4804 11228 4856 11280
rect 8300 11271 8352 11280
rect 8300 11237 8309 11271
rect 8309 11237 8343 11271
rect 8343 11237 8352 11271
rect 8300 11228 8352 11237
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 3056 11160 3108 11212
rect 3148 11024 3200 11076
rect 5448 11160 5500 11212
rect 9772 11296 9824 11348
rect 10232 11339 10284 11348
rect 10232 11305 10249 11339
rect 10249 11305 10284 11339
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 8852 11203 8904 11212
rect 8852 11169 8861 11203
rect 8861 11169 8895 11203
rect 8895 11169 8904 11203
rect 8852 11160 8904 11169
rect 9496 11228 9548 11280
rect 10232 11296 10284 11305
rect 10416 11271 10468 11280
rect 10416 11237 10425 11271
rect 10425 11237 10459 11271
rect 10459 11237 10468 11271
rect 10416 11228 10468 11237
rect 13084 11228 13136 11280
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 10324 11160 10376 11212
rect 11336 11160 11388 11212
rect 12624 11203 12676 11212
rect 12624 11169 12633 11203
rect 12633 11169 12667 11203
rect 12667 11169 12676 11203
rect 12624 11160 12676 11169
rect 13360 11160 13412 11212
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 15292 11228 15344 11280
rect 15936 11296 15988 11348
rect 16028 11296 16080 11348
rect 16488 11296 16540 11348
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 11428 11092 11480 11144
rect 14464 11092 14516 11144
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 3332 10956 3384 11008
rect 4896 10956 4948 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 10140 11024 10192 11076
rect 13820 11024 13872 11076
rect 15108 11203 15160 11212
rect 15108 11169 15117 11203
rect 15117 11169 15151 11203
rect 15151 11169 15160 11203
rect 15476 11203 15528 11212
rect 15108 11160 15160 11169
rect 15476 11169 15485 11203
rect 15485 11169 15519 11203
rect 15519 11169 15528 11203
rect 15476 11160 15528 11169
rect 15660 11203 15712 11212
rect 15660 11169 15669 11203
rect 15669 11169 15703 11203
rect 15703 11169 15712 11203
rect 15660 11160 15712 11169
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 16028 11160 16080 11212
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 16672 11160 16724 11212
rect 16856 11203 16908 11212
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 17224 11160 17276 11212
rect 16396 11024 16448 11076
rect 14464 10999 14516 11008
rect 14464 10965 14473 10999
rect 14473 10965 14507 10999
rect 14507 10965 14516 10999
rect 14464 10956 14516 10965
rect 15108 10956 15160 11008
rect 15292 10956 15344 11008
rect 15568 10956 15620 11008
rect 2755 10854 2807 10906
rect 2819 10854 2871 10906
rect 2883 10854 2935 10906
rect 2947 10854 2999 10906
rect 3011 10854 3063 10906
rect 7470 10854 7522 10906
rect 7534 10854 7586 10906
rect 7598 10854 7650 10906
rect 7662 10854 7714 10906
rect 7726 10854 7778 10906
rect 12185 10854 12237 10906
rect 12249 10854 12301 10906
rect 12313 10854 12365 10906
rect 12377 10854 12429 10906
rect 12441 10854 12493 10906
rect 16900 10854 16952 10906
rect 16964 10854 17016 10906
rect 17028 10854 17080 10906
rect 17092 10854 17144 10906
rect 17156 10854 17208 10906
rect 3148 10752 3200 10804
rect 9496 10752 9548 10804
rect 13268 10752 13320 10804
rect 14464 10795 14516 10804
rect 14464 10761 14473 10795
rect 14473 10761 14507 10795
rect 14507 10761 14516 10795
rect 14464 10752 14516 10761
rect 14740 10752 14792 10804
rect 15476 10752 15528 10804
rect 15844 10752 15896 10804
rect 9680 10684 9732 10736
rect 11244 10684 11296 10736
rect 13452 10684 13504 10736
rect 1768 10548 1820 10600
rect 1860 10480 1912 10532
rect 7380 10548 7432 10600
rect 8024 10616 8076 10668
rect 11336 10659 11388 10668
rect 11336 10625 11345 10659
rect 11345 10625 11379 10659
rect 11379 10625 11388 10659
rect 11336 10616 11388 10625
rect 12808 10616 12860 10668
rect 14188 10684 14240 10736
rect 15016 10684 15068 10736
rect 15292 10684 15344 10736
rect 7932 10548 7984 10600
rect 8392 10591 8444 10600
rect 8392 10557 8401 10591
rect 8401 10557 8435 10591
rect 8435 10557 8444 10591
rect 8392 10548 8444 10557
rect 9036 10548 9088 10600
rect 11428 10591 11480 10600
rect 11428 10557 11437 10591
rect 11437 10557 11471 10591
rect 11471 10557 11480 10591
rect 11428 10548 11480 10557
rect 12624 10548 12676 10600
rect 13636 10548 13688 10600
rect 13360 10480 13412 10532
rect 14188 10548 14240 10600
rect 15660 10616 15712 10668
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 15108 10591 15160 10600
rect 15108 10557 15117 10591
rect 15117 10557 15151 10591
rect 15151 10557 15160 10591
rect 15108 10548 15160 10557
rect 15844 10548 15896 10600
rect 16304 10616 16356 10668
rect 16396 10616 16448 10668
rect 17224 10684 17276 10736
rect 16764 10548 16816 10600
rect 17500 10548 17552 10600
rect 8300 10412 8352 10464
rect 13544 10455 13596 10464
rect 13544 10421 13553 10455
rect 13553 10421 13587 10455
rect 13587 10421 13596 10455
rect 13544 10412 13596 10421
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 14004 10412 14056 10464
rect 14372 10412 14424 10464
rect 15016 10412 15068 10464
rect 15200 10412 15252 10464
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 16028 10455 16080 10464
rect 16028 10421 16037 10455
rect 16037 10421 16071 10455
rect 16071 10421 16080 10455
rect 16028 10412 16080 10421
rect 16488 10412 16540 10464
rect 17868 10412 17920 10464
rect 5112 10310 5164 10362
rect 5176 10310 5228 10362
rect 5240 10310 5292 10362
rect 5304 10310 5356 10362
rect 5368 10310 5420 10362
rect 9827 10310 9879 10362
rect 9891 10310 9943 10362
rect 9955 10310 10007 10362
rect 10019 10310 10071 10362
rect 10083 10310 10135 10362
rect 14542 10310 14594 10362
rect 14606 10310 14658 10362
rect 14670 10310 14722 10362
rect 14734 10310 14786 10362
rect 14798 10310 14850 10362
rect 19257 10310 19309 10362
rect 19321 10310 19373 10362
rect 19385 10310 19437 10362
rect 19449 10310 19501 10362
rect 19513 10310 19565 10362
rect 10692 10208 10744 10260
rect 13636 10208 13688 10260
rect 14188 10251 14240 10260
rect 14188 10217 14197 10251
rect 14197 10217 14231 10251
rect 14231 10217 14240 10251
rect 14188 10208 14240 10217
rect 15200 10208 15252 10260
rect 15384 10208 15436 10260
rect 17868 10251 17920 10260
rect 17868 10217 17877 10251
rect 17877 10217 17911 10251
rect 17911 10217 17920 10251
rect 17868 10208 17920 10217
rect 7012 10072 7064 10124
rect 7380 10115 7432 10124
rect 7380 10081 7389 10115
rect 7389 10081 7423 10115
rect 7423 10081 7432 10115
rect 7380 10072 7432 10081
rect 8208 10072 8260 10124
rect 9496 10072 9548 10124
rect 9956 10072 10008 10124
rect 10140 10072 10192 10124
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 12624 10072 12676 10124
rect 13176 10115 13228 10124
rect 13176 10081 13185 10115
rect 13185 10081 13219 10115
rect 13219 10081 13228 10115
rect 13176 10072 13228 10081
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13912 10140 13964 10192
rect 15752 10140 15804 10192
rect 16028 10140 16080 10192
rect 13636 10115 13688 10124
rect 13636 10081 13645 10115
rect 13645 10081 13679 10115
rect 13679 10081 13688 10115
rect 13636 10072 13688 10081
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10324 10004 10376 10056
rect 10140 9936 10192 9988
rect 12900 9979 12952 9988
rect 12900 9945 12909 9979
rect 12909 9945 12943 9979
rect 12943 9945 12952 9979
rect 14004 10047 14056 10056
rect 14004 10013 14013 10047
rect 14013 10013 14047 10047
rect 14047 10013 14056 10047
rect 14004 10004 14056 10013
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 14648 10072 14700 10124
rect 16212 10072 16264 10124
rect 17316 10072 17368 10124
rect 12900 9936 12952 9945
rect 7380 9868 7432 9920
rect 9496 9868 9548 9920
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 13268 9868 13320 9920
rect 16120 10004 16172 10056
rect 14740 9979 14792 9988
rect 14740 9945 14749 9979
rect 14749 9945 14783 9979
rect 14783 9945 14792 9979
rect 14740 9936 14792 9945
rect 16580 9936 16632 9988
rect 16304 9868 16356 9920
rect 17316 9868 17368 9920
rect 17868 9868 17920 9920
rect 2755 9766 2807 9818
rect 2819 9766 2871 9818
rect 2883 9766 2935 9818
rect 2947 9766 2999 9818
rect 3011 9766 3063 9818
rect 7470 9766 7522 9818
rect 7534 9766 7586 9818
rect 7598 9766 7650 9818
rect 7662 9766 7714 9818
rect 7726 9766 7778 9818
rect 12185 9766 12237 9818
rect 12249 9766 12301 9818
rect 12313 9766 12365 9818
rect 12377 9766 12429 9818
rect 12441 9766 12493 9818
rect 16900 9766 16952 9818
rect 16964 9766 17016 9818
rect 17028 9766 17080 9818
rect 17092 9766 17144 9818
rect 17156 9766 17208 9818
rect 9956 9664 10008 9716
rect 10232 9664 10284 9716
rect 12624 9664 12676 9716
rect 8392 9528 8444 9580
rect 12992 9596 13044 9648
rect 14096 9707 14148 9716
rect 14096 9673 14105 9707
rect 14105 9673 14139 9707
rect 14139 9673 14148 9707
rect 14096 9664 14148 9673
rect 14372 9664 14424 9716
rect 15200 9664 15252 9716
rect 16488 9664 16540 9716
rect 16672 9596 16724 9648
rect 9772 9460 9824 9512
rect 7656 9435 7708 9444
rect 7656 9401 7674 9435
rect 7674 9401 7708 9435
rect 7656 9392 7708 9401
rect 6184 9324 6236 9376
rect 7472 9324 7524 9376
rect 9496 9324 9548 9376
rect 9956 9503 10008 9512
rect 9956 9469 9965 9503
rect 9965 9469 9999 9503
rect 9999 9469 10008 9503
rect 9956 9460 10008 9469
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10140 9460 10192 9512
rect 11428 9528 11480 9580
rect 12716 9528 12768 9580
rect 13176 9528 13228 9580
rect 11244 9460 11296 9512
rect 10416 9324 10468 9376
rect 11888 9324 11940 9376
rect 13728 9503 13780 9512
rect 13728 9469 13737 9503
rect 13737 9469 13771 9503
rect 13771 9469 13780 9503
rect 13728 9460 13780 9469
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 14464 9528 14516 9580
rect 15384 9528 15436 9580
rect 15200 9460 15252 9512
rect 15752 9460 15804 9512
rect 17316 9528 17368 9580
rect 16304 9503 16356 9512
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 16672 9460 16724 9512
rect 16212 9392 16264 9444
rect 15200 9324 15252 9376
rect 15292 9324 15344 9376
rect 5112 9222 5164 9274
rect 5176 9222 5228 9274
rect 5240 9222 5292 9274
rect 5304 9222 5356 9274
rect 5368 9222 5420 9274
rect 9827 9222 9879 9274
rect 9891 9222 9943 9274
rect 9955 9222 10007 9274
rect 10019 9222 10071 9274
rect 10083 9222 10135 9274
rect 14542 9222 14594 9274
rect 14606 9222 14658 9274
rect 14670 9222 14722 9274
rect 14734 9222 14786 9274
rect 14798 9222 14850 9274
rect 19257 9222 19309 9274
rect 19321 9222 19373 9274
rect 19385 9222 19437 9274
rect 19449 9222 19501 9274
rect 19513 9222 19565 9274
rect 7380 9120 7432 9172
rect 11520 9120 11572 9172
rect 12900 9120 12952 9172
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 8944 9052 8996 9104
rect 7472 8984 7524 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 10232 8984 10284 9036
rect 17224 9120 17276 9172
rect 10416 8916 10468 8968
rect 11520 8984 11572 9036
rect 11796 9027 11848 9036
rect 11796 8993 11805 9027
rect 11805 8993 11839 9027
rect 11839 8993 11848 9027
rect 11796 8984 11848 8993
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 7656 8891 7708 8900
rect 7656 8857 7665 8891
rect 7665 8857 7699 8891
rect 7699 8857 7708 8891
rect 7656 8848 7708 8857
rect 12532 8984 12584 9036
rect 13084 9027 13136 9036
rect 13084 8993 13093 9027
rect 13093 8993 13127 9027
rect 13127 8993 13136 9027
rect 13084 8984 13136 8993
rect 13176 9027 13228 9036
rect 13176 8993 13185 9027
rect 13185 8993 13219 9027
rect 13219 8993 13228 9027
rect 13176 8984 13228 8993
rect 13728 8984 13780 9036
rect 15660 9027 15712 9036
rect 15660 8993 15669 9027
rect 15669 8993 15703 9027
rect 15703 8993 15712 9027
rect 15660 8984 15712 8993
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 17316 8984 17368 9036
rect 18328 8984 18380 9036
rect 12716 8916 12768 8968
rect 15844 8916 15896 8968
rect 12624 8848 12676 8900
rect 15016 8848 15068 8900
rect 17224 8916 17276 8968
rect 17408 8959 17460 8968
rect 17408 8925 17417 8959
rect 17417 8925 17451 8959
rect 17451 8925 17460 8959
rect 17408 8916 17460 8925
rect 8852 8823 8904 8832
rect 8852 8789 8861 8823
rect 8861 8789 8895 8823
rect 8895 8789 8904 8823
rect 8852 8780 8904 8789
rect 10324 8780 10376 8832
rect 15384 8780 15436 8832
rect 16120 8780 16172 8832
rect 2755 8678 2807 8730
rect 2819 8678 2871 8730
rect 2883 8678 2935 8730
rect 2947 8678 2999 8730
rect 3011 8678 3063 8730
rect 7470 8678 7522 8730
rect 7534 8678 7586 8730
rect 7598 8678 7650 8730
rect 7662 8678 7714 8730
rect 7726 8678 7778 8730
rect 12185 8678 12237 8730
rect 12249 8678 12301 8730
rect 12313 8678 12365 8730
rect 12377 8678 12429 8730
rect 12441 8678 12493 8730
rect 16900 8678 16952 8730
rect 16964 8678 17016 8730
rect 17028 8678 17080 8730
rect 17092 8678 17144 8730
rect 17156 8678 17208 8730
rect 11796 8576 11848 8628
rect 13176 8576 13228 8628
rect 14096 8576 14148 8628
rect 16764 8576 16816 8628
rect 18328 8619 18380 8628
rect 8668 8508 8720 8560
rect 13268 8440 13320 8492
rect 8392 8372 8444 8424
rect 12532 8372 12584 8424
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 13820 8372 13872 8424
rect 15016 8508 15068 8560
rect 8852 8304 8904 8356
rect 9772 8304 9824 8356
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 14924 8440 14976 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16672 8440 16724 8492
rect 14096 8279 14148 8288
rect 14096 8245 14105 8279
rect 14105 8245 14139 8279
rect 14139 8245 14148 8279
rect 14096 8236 14148 8245
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 15660 8372 15712 8424
rect 15752 8415 15804 8424
rect 15752 8381 15761 8415
rect 15761 8381 15795 8415
rect 15795 8381 15804 8415
rect 15752 8372 15804 8381
rect 15844 8415 15896 8424
rect 15844 8381 15853 8415
rect 15853 8381 15887 8415
rect 15887 8381 15896 8415
rect 15844 8372 15896 8381
rect 16028 8415 16080 8424
rect 16028 8381 16037 8415
rect 16037 8381 16071 8415
rect 16071 8381 16080 8415
rect 16028 8372 16080 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 16580 8372 16632 8424
rect 16856 8372 16908 8424
rect 17408 8440 17460 8492
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 17960 8440 18012 8492
rect 16396 8304 16448 8356
rect 15476 8236 15528 8288
rect 16304 8236 16356 8288
rect 16764 8236 16816 8288
rect 17868 8236 17920 8288
rect 18052 8304 18104 8356
rect 5112 8134 5164 8186
rect 5176 8134 5228 8186
rect 5240 8134 5292 8186
rect 5304 8134 5356 8186
rect 5368 8134 5420 8186
rect 9827 8134 9879 8186
rect 9891 8134 9943 8186
rect 9955 8134 10007 8186
rect 10019 8134 10071 8186
rect 10083 8134 10135 8186
rect 14542 8134 14594 8186
rect 14606 8134 14658 8186
rect 14670 8134 14722 8186
rect 14734 8134 14786 8186
rect 14798 8134 14850 8186
rect 19257 8134 19309 8186
rect 19321 8134 19373 8186
rect 19385 8134 19437 8186
rect 19449 8134 19501 8186
rect 19513 8134 19565 8186
rect 9864 8032 9916 8084
rect 10324 8032 10376 8084
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 12716 8032 12768 8084
rect 9496 7964 9548 8016
rect 12532 7964 12584 8016
rect 13544 8032 13596 8084
rect 15752 8032 15804 8084
rect 15936 8032 15988 8084
rect 16304 8032 16356 8084
rect 12900 7896 12952 7948
rect 13176 7939 13228 7948
rect 13176 7905 13185 7939
rect 13185 7905 13219 7939
rect 13219 7905 13228 7939
rect 13176 7896 13228 7905
rect 13544 7896 13596 7948
rect 15016 7964 15068 8016
rect 15476 7896 15528 7948
rect 16396 7939 16448 7948
rect 16396 7905 16405 7939
rect 16405 7905 16439 7939
rect 16439 7905 16448 7939
rect 16396 7896 16448 7905
rect 14832 7828 14884 7880
rect 17500 7964 17552 8016
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 14924 7760 14976 7812
rect 15200 7760 15252 7812
rect 16580 7760 16632 7812
rect 16856 7760 16908 7812
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 12900 7692 12952 7744
rect 15016 7692 15068 7744
rect 15108 7692 15160 7744
rect 17868 7896 17920 7948
rect 2755 7590 2807 7642
rect 2819 7590 2871 7642
rect 2883 7590 2935 7642
rect 2947 7590 2999 7642
rect 3011 7590 3063 7642
rect 7470 7590 7522 7642
rect 7534 7590 7586 7642
rect 7598 7590 7650 7642
rect 7662 7590 7714 7642
rect 7726 7590 7778 7642
rect 12185 7590 12237 7642
rect 12249 7590 12301 7642
rect 12313 7590 12365 7642
rect 12377 7590 12429 7642
rect 12441 7590 12493 7642
rect 16900 7590 16952 7642
rect 16964 7590 17016 7642
rect 17028 7590 17080 7642
rect 17092 7590 17144 7642
rect 17156 7590 17208 7642
rect 13912 7488 13964 7540
rect 14832 7488 14884 7540
rect 15568 7488 15620 7540
rect 16764 7488 16816 7540
rect 8392 7420 8444 7472
rect 8484 7284 8536 7336
rect 8944 7284 8996 7336
rect 9496 7284 9548 7336
rect 6552 7259 6604 7268
rect 6552 7225 6561 7259
rect 6561 7225 6595 7259
rect 6595 7225 6604 7259
rect 6552 7216 6604 7225
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 8300 7148 8352 7200
rect 10324 7148 10376 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 12808 7420 12860 7472
rect 13176 7420 13228 7472
rect 14280 7420 14332 7472
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12624 7284 12676 7336
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 12992 7284 13044 7336
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 13176 7327 13228 7336
rect 13176 7293 13185 7327
rect 13185 7293 13219 7327
rect 13219 7293 13228 7327
rect 13176 7284 13228 7293
rect 12072 7259 12124 7268
rect 12072 7225 12081 7259
rect 12081 7225 12115 7259
rect 12115 7225 12124 7259
rect 12072 7216 12124 7225
rect 12164 7259 12216 7268
rect 12164 7225 12173 7259
rect 12173 7225 12207 7259
rect 12207 7225 12216 7259
rect 12164 7216 12216 7225
rect 12808 7259 12860 7268
rect 12808 7225 12817 7259
rect 12817 7225 12851 7259
rect 12851 7225 12860 7259
rect 12808 7216 12860 7225
rect 13544 7352 13596 7404
rect 13452 7216 13504 7268
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 14464 7352 14516 7404
rect 14832 7284 14884 7336
rect 15108 7352 15160 7404
rect 15016 7327 15068 7336
rect 15016 7293 15025 7327
rect 15025 7293 15059 7327
rect 15059 7293 15068 7327
rect 15016 7284 15068 7293
rect 16488 7420 16540 7472
rect 14096 7148 14148 7200
rect 14372 7148 14424 7200
rect 14464 7191 14516 7200
rect 14464 7157 14473 7191
rect 14473 7157 14507 7191
rect 14507 7157 14516 7191
rect 14464 7148 14516 7157
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 17224 7352 17276 7404
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 16396 7148 16448 7200
rect 5112 7046 5164 7098
rect 5176 7046 5228 7098
rect 5240 7046 5292 7098
rect 5304 7046 5356 7098
rect 5368 7046 5420 7098
rect 9827 7046 9879 7098
rect 9891 7046 9943 7098
rect 9955 7046 10007 7098
rect 10019 7046 10071 7098
rect 10083 7046 10135 7098
rect 14542 7046 14594 7098
rect 14606 7046 14658 7098
rect 14670 7046 14722 7098
rect 14734 7046 14786 7098
rect 14798 7046 14850 7098
rect 19257 7046 19309 7098
rect 19321 7046 19373 7098
rect 19385 7046 19437 7098
rect 19449 7046 19501 7098
rect 19513 7046 19565 7098
rect 9680 6944 9732 6996
rect 12072 6944 12124 6996
rect 12624 6987 12676 6996
rect 12624 6953 12633 6987
rect 12633 6953 12667 6987
rect 12667 6953 12676 6987
rect 12624 6944 12676 6953
rect 13084 6944 13136 6996
rect 13452 6944 13504 6996
rect 13820 6944 13872 6996
rect 14280 6944 14332 6996
rect 8944 6876 8996 6928
rect 9496 6876 9548 6928
rect 11520 6876 11572 6928
rect 8576 6808 8628 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11152 6808 11204 6860
rect 11336 6808 11388 6860
rect 12532 6808 12584 6860
rect 12716 6851 12768 6860
rect 12716 6817 12725 6851
rect 12725 6817 12759 6851
rect 12759 6817 12768 6851
rect 12716 6808 12768 6817
rect 11796 6740 11848 6792
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 13820 6808 13872 6860
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 14280 6851 14332 6860
rect 14280 6817 14289 6851
rect 14289 6817 14323 6851
rect 14323 6817 14332 6851
rect 14280 6808 14332 6817
rect 14464 6808 14516 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15200 6851 15252 6860
rect 15200 6817 15209 6851
rect 15209 6817 15243 6851
rect 15243 6817 15252 6851
rect 15200 6808 15252 6817
rect 15292 6851 15344 6860
rect 15292 6817 15301 6851
rect 15301 6817 15335 6851
rect 15335 6817 15344 6851
rect 15292 6808 15344 6817
rect 15568 6876 15620 6928
rect 15660 6876 15712 6928
rect 16488 6808 16540 6860
rect 16028 6740 16080 6792
rect 16396 6783 16448 6792
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 9588 6604 9640 6656
rect 9956 6604 10008 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 15200 6672 15252 6724
rect 2755 6502 2807 6554
rect 2819 6502 2871 6554
rect 2883 6502 2935 6554
rect 2947 6502 2999 6554
rect 3011 6502 3063 6554
rect 7470 6502 7522 6554
rect 7534 6502 7586 6554
rect 7598 6502 7650 6554
rect 7662 6502 7714 6554
rect 7726 6502 7778 6554
rect 12185 6502 12237 6554
rect 12249 6502 12301 6554
rect 12313 6502 12365 6554
rect 12377 6502 12429 6554
rect 12441 6502 12493 6554
rect 16900 6502 16952 6554
rect 16964 6502 17016 6554
rect 17028 6502 17080 6554
rect 17092 6502 17144 6554
rect 17156 6502 17208 6554
rect 8944 6400 8996 6452
rect 8392 6196 8444 6248
rect 9312 6196 9364 6248
rect 9956 6239 10008 6248
rect 9956 6205 9965 6239
rect 9965 6205 9999 6239
rect 9999 6205 10008 6239
rect 9956 6196 10008 6205
rect 12532 6400 12584 6452
rect 14556 6400 14608 6452
rect 10232 6375 10284 6384
rect 10232 6341 10241 6375
rect 10241 6341 10275 6375
rect 10275 6341 10284 6375
rect 10232 6332 10284 6341
rect 11520 6332 11572 6384
rect 9588 6171 9640 6180
rect 9588 6137 9606 6171
rect 9606 6137 9640 6171
rect 10324 6239 10376 6248
rect 10324 6205 10333 6239
rect 10333 6205 10367 6239
rect 10367 6205 10376 6239
rect 10324 6196 10376 6205
rect 10692 6196 10744 6248
rect 9588 6128 9640 6137
rect 11336 6128 11388 6180
rect 8484 6103 8536 6112
rect 8484 6069 8493 6103
rect 8493 6069 8527 6103
rect 8527 6069 8536 6103
rect 8484 6060 8536 6069
rect 9404 6060 9456 6112
rect 5112 5958 5164 6010
rect 5176 5958 5228 6010
rect 5240 5958 5292 6010
rect 5304 5958 5356 6010
rect 5368 5958 5420 6010
rect 9827 5958 9879 6010
rect 9891 5958 9943 6010
rect 9955 5958 10007 6010
rect 10019 5958 10071 6010
rect 10083 5958 10135 6010
rect 14542 5958 14594 6010
rect 14606 5958 14658 6010
rect 14670 5958 14722 6010
rect 14734 5958 14786 6010
rect 14798 5958 14850 6010
rect 19257 5958 19309 6010
rect 19321 5958 19373 6010
rect 19385 5958 19437 6010
rect 19449 5958 19501 6010
rect 19513 5958 19565 6010
rect 9312 5763 9364 5772
rect 9312 5729 9321 5763
rect 9321 5729 9355 5763
rect 9355 5729 9364 5763
rect 9312 5720 9364 5729
rect 10140 5720 10192 5772
rect 11060 5720 11112 5772
rect 11520 5720 11572 5772
rect 16580 5788 16632 5840
rect 11152 5516 11204 5568
rect 16120 5516 16172 5568
rect 18604 5516 18656 5568
rect 2755 5414 2807 5466
rect 2819 5414 2871 5466
rect 2883 5414 2935 5466
rect 2947 5414 2999 5466
rect 3011 5414 3063 5466
rect 7470 5414 7522 5466
rect 7534 5414 7586 5466
rect 7598 5414 7650 5466
rect 7662 5414 7714 5466
rect 7726 5414 7778 5466
rect 12185 5414 12237 5466
rect 12249 5414 12301 5466
rect 12313 5414 12365 5466
rect 12377 5414 12429 5466
rect 12441 5414 12493 5466
rect 16900 5414 16952 5466
rect 16964 5414 17016 5466
rect 17028 5414 17080 5466
rect 17092 5414 17144 5466
rect 17156 5414 17208 5466
rect 11060 5176 11112 5228
rect 11244 5108 11296 5160
rect 13636 4972 13688 5024
rect 5112 4870 5164 4922
rect 5176 4870 5228 4922
rect 5240 4870 5292 4922
rect 5304 4870 5356 4922
rect 5368 4870 5420 4922
rect 9827 4870 9879 4922
rect 9891 4870 9943 4922
rect 9955 4870 10007 4922
rect 10019 4870 10071 4922
rect 10083 4870 10135 4922
rect 14542 4870 14594 4922
rect 14606 4870 14658 4922
rect 14670 4870 14722 4922
rect 14734 4870 14786 4922
rect 14798 4870 14850 4922
rect 19257 4870 19309 4922
rect 19321 4870 19373 4922
rect 19385 4870 19437 4922
rect 19449 4870 19501 4922
rect 19513 4870 19565 4922
rect 2755 4326 2807 4378
rect 2819 4326 2871 4378
rect 2883 4326 2935 4378
rect 2947 4326 2999 4378
rect 3011 4326 3063 4378
rect 7470 4326 7522 4378
rect 7534 4326 7586 4378
rect 7598 4326 7650 4378
rect 7662 4326 7714 4378
rect 7726 4326 7778 4378
rect 12185 4326 12237 4378
rect 12249 4326 12301 4378
rect 12313 4326 12365 4378
rect 12377 4326 12429 4378
rect 12441 4326 12493 4378
rect 16900 4326 16952 4378
rect 16964 4326 17016 4378
rect 17028 4326 17080 4378
rect 17092 4326 17144 4378
rect 17156 4326 17208 4378
rect 3700 4088 3752 4140
rect 8484 4088 8536 4140
rect 5112 3782 5164 3834
rect 5176 3782 5228 3834
rect 5240 3782 5292 3834
rect 5304 3782 5356 3834
rect 5368 3782 5420 3834
rect 9827 3782 9879 3834
rect 9891 3782 9943 3834
rect 9955 3782 10007 3834
rect 10019 3782 10071 3834
rect 10083 3782 10135 3834
rect 14542 3782 14594 3834
rect 14606 3782 14658 3834
rect 14670 3782 14722 3834
rect 14734 3782 14786 3834
rect 14798 3782 14850 3834
rect 19257 3782 19309 3834
rect 19321 3782 19373 3834
rect 19385 3782 19437 3834
rect 19449 3782 19501 3834
rect 19513 3782 19565 3834
rect 1216 3476 1268 3528
rect 6552 3476 6604 3528
rect 2755 3238 2807 3290
rect 2819 3238 2871 3290
rect 2883 3238 2935 3290
rect 2947 3238 2999 3290
rect 3011 3238 3063 3290
rect 7470 3238 7522 3290
rect 7534 3238 7586 3290
rect 7598 3238 7650 3290
rect 7662 3238 7714 3290
rect 7726 3238 7778 3290
rect 12185 3238 12237 3290
rect 12249 3238 12301 3290
rect 12313 3238 12365 3290
rect 12377 3238 12429 3290
rect 12441 3238 12493 3290
rect 16900 3238 16952 3290
rect 16964 3238 17016 3290
rect 17028 3238 17080 3290
rect 17092 3238 17144 3290
rect 17156 3238 17208 3290
rect 5112 2694 5164 2746
rect 5176 2694 5228 2746
rect 5240 2694 5292 2746
rect 5304 2694 5356 2746
rect 5368 2694 5420 2746
rect 9827 2694 9879 2746
rect 9891 2694 9943 2746
rect 9955 2694 10007 2746
rect 10019 2694 10071 2746
rect 10083 2694 10135 2746
rect 14542 2694 14594 2746
rect 14606 2694 14658 2746
rect 14670 2694 14722 2746
rect 14734 2694 14786 2746
rect 14798 2694 14850 2746
rect 19257 2694 19309 2746
rect 19321 2694 19373 2746
rect 19385 2694 19437 2746
rect 19449 2694 19501 2746
rect 19513 2694 19565 2746
rect 2755 2150 2807 2202
rect 2819 2150 2871 2202
rect 2883 2150 2935 2202
rect 2947 2150 2999 2202
rect 3011 2150 3063 2202
rect 7470 2150 7522 2202
rect 7534 2150 7586 2202
rect 7598 2150 7650 2202
rect 7662 2150 7714 2202
rect 7726 2150 7778 2202
rect 12185 2150 12237 2202
rect 12249 2150 12301 2202
rect 12313 2150 12365 2202
rect 12377 2150 12429 2202
rect 12441 2150 12493 2202
rect 16900 2150 16952 2202
rect 16964 2150 17016 2202
rect 17028 2150 17080 2202
rect 17092 2150 17144 2202
rect 17156 2150 17208 2202
rect 5112 1606 5164 1658
rect 5176 1606 5228 1658
rect 5240 1606 5292 1658
rect 5304 1606 5356 1658
rect 5368 1606 5420 1658
rect 9827 1606 9879 1658
rect 9891 1606 9943 1658
rect 9955 1606 10007 1658
rect 10019 1606 10071 1658
rect 10083 1606 10135 1658
rect 14542 1606 14594 1658
rect 14606 1606 14658 1658
rect 14670 1606 14722 1658
rect 14734 1606 14786 1658
rect 14798 1606 14850 1658
rect 19257 1606 19309 1658
rect 19321 1606 19373 1658
rect 19385 1606 19437 1658
rect 19449 1606 19501 1658
rect 19513 1606 19565 1658
rect 2755 1062 2807 1114
rect 2819 1062 2871 1114
rect 2883 1062 2935 1114
rect 2947 1062 2999 1114
rect 3011 1062 3063 1114
rect 7470 1062 7522 1114
rect 7534 1062 7586 1114
rect 7598 1062 7650 1114
rect 7662 1062 7714 1114
rect 7726 1062 7778 1114
rect 12185 1062 12237 1114
rect 12249 1062 12301 1114
rect 12313 1062 12365 1114
rect 12377 1062 12429 1114
rect 12441 1062 12493 1114
rect 16900 1062 16952 1114
rect 16964 1062 17016 1114
rect 17028 1062 17080 1114
rect 17092 1062 17144 1114
rect 17156 1062 17208 1114
rect 5112 518 5164 570
rect 5176 518 5228 570
rect 5240 518 5292 570
rect 5304 518 5356 570
rect 5368 518 5420 570
rect 9827 518 9879 570
rect 9891 518 9943 570
rect 9955 518 10007 570
rect 10019 518 10071 570
rect 10083 518 10135 570
rect 14542 518 14594 570
rect 14606 518 14658 570
rect 14670 518 14722 570
rect 14734 518 14786 570
rect 14798 518 14850 570
rect 19257 518 19309 570
rect 19321 518 19373 570
rect 19385 518 19437 570
rect 19449 518 19501 570
rect 19513 518 19565 570
<< metal2 >>
rect 846 19600 902 20000
rect 2502 19600 2558 20000
rect 4158 19600 4214 20000
rect 5814 19600 5870 20000
rect 7470 19600 7526 20000
rect 9126 19600 9182 20000
rect 10782 19600 10838 20000
rect 12438 19600 12494 20000
rect 14094 19600 14150 20000
rect 15750 19600 15806 20000
rect 17406 19600 17462 20000
rect 19062 19600 19118 20000
rect 860 18834 888 19600
rect 2516 18834 2544 19600
rect 4172 18834 4200 19600
rect 5112 19068 5420 19077
rect 5112 19066 5118 19068
rect 5174 19066 5198 19068
rect 5254 19066 5278 19068
rect 5334 19066 5358 19068
rect 5414 19066 5420 19068
rect 5174 19014 5176 19066
rect 5356 19014 5358 19066
rect 5112 19012 5118 19014
rect 5174 19012 5198 19014
rect 5254 19012 5278 19014
rect 5334 19012 5358 19014
rect 5414 19012 5420 19014
rect 5112 19003 5420 19012
rect 5828 18834 5856 19600
rect 7484 18834 7512 19600
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 848 18828 900 18834
rect 848 18770 900 18776
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 5816 18828 5868 18834
rect 5816 18770 5868 18776
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 2755 18524 3063 18533
rect 2755 18522 2761 18524
rect 2817 18522 2841 18524
rect 2897 18522 2921 18524
rect 2977 18522 3001 18524
rect 3057 18522 3063 18524
rect 2817 18470 2819 18522
rect 2999 18470 3001 18522
rect 2755 18468 2761 18470
rect 2817 18468 2841 18470
rect 2897 18468 2921 18470
rect 2977 18468 3001 18470
rect 3057 18468 3063 18470
rect 2755 18459 3063 18468
rect 3608 18216 3660 18222
rect 3608 18158 3660 18164
rect 3792 18216 3844 18222
rect 3792 18158 3844 18164
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 848 17672 900 17678
rect 848 17614 900 17620
rect 860 15026 888 17614
rect 2056 17134 2084 17818
rect 3344 17746 3372 18022
rect 2320 17740 2372 17746
rect 2320 17682 2372 17688
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1308 15904 1360 15910
rect 1308 15846 1360 15852
rect 1320 15366 1348 15846
rect 1780 15638 1808 16050
rect 2056 16028 2084 17070
rect 2148 16182 2176 17070
rect 2332 16794 2360 17682
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 2755 17436 3063 17445
rect 2755 17434 2761 17436
rect 2817 17434 2841 17436
rect 2897 17434 2921 17436
rect 2977 17434 3001 17436
rect 3057 17434 3063 17436
rect 2817 17382 2819 17434
rect 2999 17382 3001 17434
rect 2755 17380 2761 17382
rect 2817 17380 2841 17382
rect 2897 17380 2921 17382
rect 2977 17380 3001 17382
rect 3057 17380 3063 17382
rect 2755 17371 3063 17380
rect 3252 17134 3280 17478
rect 3620 17338 3648 18158
rect 3804 17814 3832 18158
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 3792 17808 3844 17814
rect 3792 17750 3844 17756
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2516 16658 2544 16934
rect 3252 16658 3280 17070
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2755 16348 3063 16357
rect 2755 16346 2761 16348
rect 2817 16346 2841 16348
rect 2897 16346 2921 16348
rect 2977 16346 3001 16348
rect 3057 16346 3063 16348
rect 2817 16294 2819 16346
rect 2999 16294 3001 16346
rect 2755 16292 2761 16294
rect 2817 16292 2841 16294
rect 2897 16292 2921 16294
rect 2977 16292 3001 16294
rect 3057 16292 3063 16294
rect 2755 16283 3063 16292
rect 2136 16176 2188 16182
rect 2136 16118 2188 16124
rect 2136 16040 2188 16046
rect 2056 16000 2136 16028
rect 2136 15982 2188 15988
rect 2412 16040 2464 16046
rect 2412 15982 2464 15988
rect 2148 15706 2176 15982
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 1768 15632 1820 15638
rect 1768 15574 1820 15580
rect 1032 15360 1084 15366
rect 1032 15302 1084 15308
rect 1308 15360 1360 15366
rect 1308 15302 1360 15308
rect 848 15020 900 15026
rect 848 14962 900 14968
rect 1044 14890 1072 15302
rect 1032 14884 1084 14890
rect 1032 14826 1084 14832
rect 1780 14618 1808 15574
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1964 14346 1992 15438
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 2148 14278 2176 15642
rect 2240 15638 2268 15914
rect 2424 15706 2452 15982
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2228 15632 2280 15638
rect 2228 15574 2280 15580
rect 2240 14822 2268 15574
rect 2516 15502 2544 15914
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2596 15428 2648 15434
rect 2596 15370 2648 15376
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 14958 2360 15302
rect 2608 15042 2636 15370
rect 2755 15260 3063 15269
rect 2755 15258 2761 15260
rect 2817 15258 2841 15260
rect 2897 15258 2921 15260
rect 2977 15258 3001 15260
rect 3057 15258 3063 15260
rect 2817 15206 2819 15258
rect 2999 15206 3001 15258
rect 2755 15204 2761 15206
rect 2817 15204 2841 15206
rect 2897 15204 2921 15206
rect 2977 15204 3001 15206
rect 3057 15204 3063 15206
rect 2755 15195 3063 15204
rect 3252 15162 3280 15846
rect 3344 15706 3372 17002
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3804 15570 3832 17750
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 3976 17196 4028 17202
rect 3976 17138 4028 17144
rect 3988 16794 4016 17138
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3976 16788 4028 16794
rect 3976 16730 4028 16736
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3792 15564 3844 15570
rect 3792 15506 3844 15512
rect 3528 15162 3556 15506
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 2608 15014 2912 15042
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2884 14822 2912 15014
rect 4172 14958 4200 17070
rect 4160 14952 4212 14958
rect 4212 14912 4384 14940
rect 4160 14894 4212 14900
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 2240 14550 2268 14758
rect 2884 14550 2912 14758
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2755 14172 3063 14181
rect 2755 14170 2761 14172
rect 2817 14170 2841 14172
rect 2897 14170 2921 14172
rect 2977 14170 3001 14172
rect 3057 14170 3063 14172
rect 2817 14118 2819 14170
rect 2999 14118 3001 14170
rect 2755 14116 2761 14118
rect 2817 14116 2841 14118
rect 2897 14116 2921 14118
rect 2977 14116 3001 14118
rect 3057 14116 3063 14118
rect 2755 14107 3063 14116
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1320 13462 1348 13806
rect 1308 13456 1360 13462
rect 1308 13398 1360 13404
rect 2056 13394 2084 13806
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13530 2360 13670
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2792 13394 2820 13874
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1780 12782 1808 13126
rect 2516 12850 2544 13330
rect 2976 13190 3004 13806
rect 4080 13462 4108 14486
rect 4172 14278 4200 14758
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4356 14074 4384 14912
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14482 4568 14826
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4356 13802 4384 14010
rect 4632 13870 4660 14214
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2964 13184 3016 13190
rect 2964 13126 3016 13132
rect 2755 13084 3063 13093
rect 2755 13082 2761 13084
rect 2817 13082 2841 13084
rect 2897 13082 2921 13084
rect 2977 13082 3001 13084
rect 3057 13082 3063 13084
rect 2817 13030 2819 13082
rect 2999 13030 3001 13082
rect 2755 13028 2761 13030
rect 2817 13028 2841 13030
rect 2897 13028 2921 13030
rect 2977 13028 3001 13030
rect 3057 13028 3063 13030
rect 2755 13019 3063 13028
rect 2780 12980 2832 12986
rect 3160 12968 3188 13330
rect 4724 13326 4752 17682
rect 4908 17524 4936 17818
rect 5000 17678 5028 18022
rect 5112 17980 5420 17989
rect 5112 17978 5118 17980
rect 5174 17978 5198 17980
rect 5254 17978 5278 17980
rect 5334 17978 5358 17980
rect 5414 17978 5420 17980
rect 5174 17926 5176 17978
rect 5356 17926 5358 17978
rect 5112 17924 5118 17926
rect 5174 17924 5198 17926
rect 5254 17924 5278 17926
rect 5334 17924 5358 17926
rect 5414 17924 5420 17926
rect 5112 17915 5420 17924
rect 6472 17678 6500 18702
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 7024 18290 7052 18566
rect 7470 18524 7778 18533
rect 7470 18522 7476 18524
rect 7532 18522 7556 18524
rect 7612 18522 7636 18524
rect 7692 18522 7716 18524
rect 7772 18522 7778 18524
rect 7532 18470 7534 18522
rect 7714 18470 7716 18522
rect 7470 18468 7476 18470
rect 7532 18468 7556 18470
rect 7612 18468 7636 18470
rect 7692 18468 7716 18470
rect 7772 18468 7778 18470
rect 7470 18459 7778 18468
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 6736 18080 6788 18086
rect 6736 18022 6788 18028
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6748 17882 6776 18022
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6840 17746 6868 18022
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 5264 17536 5316 17542
rect 4908 17496 5028 17524
rect 5000 17134 5028 17496
rect 5264 17478 5316 17484
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5092 17202 5120 17274
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 5276 17134 5304 17478
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5552 17134 5580 17274
rect 5644 17134 5672 17478
rect 4988 17128 5040 17134
rect 4988 17070 5040 17076
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5000 16794 5028 17070
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5632 16992 5684 16998
rect 5632 16934 5684 16940
rect 5112 16892 5420 16901
rect 5112 16890 5118 16892
rect 5174 16890 5198 16892
rect 5254 16890 5278 16892
rect 5334 16890 5358 16892
rect 5414 16890 5420 16892
rect 5174 16838 5176 16890
rect 5356 16838 5358 16890
rect 5112 16836 5118 16838
rect 5174 16836 5198 16838
rect 5254 16836 5278 16838
rect 5334 16836 5358 16838
rect 5414 16836 5420 16838
rect 5112 16827 5420 16836
rect 4988 16788 5040 16794
rect 4988 16730 5040 16736
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 16250 5304 16526
rect 5460 16454 5488 16934
rect 5552 16658 5580 16934
rect 5644 16658 5672 16934
rect 5828 16674 5856 17070
rect 5908 17060 5960 17066
rect 5960 17020 6224 17048
rect 5908 17002 5960 17008
rect 6196 16726 6224 17020
rect 6472 16794 6500 17614
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6184 16720 6236 16726
rect 6182 16688 6184 16697
rect 6236 16688 6238 16697
rect 5828 16658 6132 16674
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5828 16652 6144 16658
rect 5828 16646 6092 16652
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5112 15804 5420 15813
rect 5112 15802 5118 15804
rect 5174 15802 5198 15804
rect 5254 15802 5278 15804
rect 5334 15802 5358 15804
rect 5414 15802 5420 15804
rect 5174 15750 5176 15802
rect 5356 15750 5358 15802
rect 5112 15748 5118 15750
rect 5174 15748 5198 15750
rect 5254 15748 5278 15750
rect 5334 15748 5358 15750
rect 5414 15748 5420 15750
rect 5112 15739 5420 15748
rect 5828 14958 5856 16646
rect 6656 16658 6684 17478
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6182 16623 6238 16632
rect 6644 16652 6696 16658
rect 6092 16594 6144 16600
rect 6644 16594 6696 16600
rect 6748 16454 6776 17274
rect 6840 17270 6868 17682
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6840 16658 6868 16730
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6288 16250 6316 16390
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 14958 6868 15846
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 4816 14006 4844 14894
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 5000 14278 5028 14758
rect 5112 14716 5420 14725
rect 5112 14714 5118 14716
rect 5174 14714 5198 14716
rect 5254 14714 5278 14716
rect 5334 14714 5358 14716
rect 5414 14714 5420 14716
rect 5174 14662 5176 14714
rect 5356 14662 5358 14714
rect 5112 14660 5118 14662
rect 5174 14660 5198 14662
rect 5254 14660 5278 14662
rect 5334 14660 5358 14662
rect 5414 14660 5420 14662
rect 5112 14651 5420 14660
rect 5828 14618 5856 14894
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5080 14544 5132 14550
rect 5080 14486 5132 14492
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 5092 13716 5120 14486
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 5184 13734 5212 14282
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13870 5396 14214
rect 5460 13870 5488 14350
rect 5552 14074 5580 14418
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5828 14006 5856 14554
rect 5816 14000 5868 14006
rect 5816 13942 5868 13948
rect 6288 13938 6316 14894
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5000 13688 5120 13716
rect 5172 13728 5224 13734
rect 5000 13512 5028 13688
rect 5172 13670 5224 13676
rect 5448 13728 5500 13734
rect 5448 13670 5500 13676
rect 5112 13628 5420 13637
rect 5112 13626 5118 13628
rect 5174 13626 5198 13628
rect 5254 13626 5278 13628
rect 5334 13626 5358 13628
rect 5414 13626 5420 13628
rect 5174 13574 5176 13626
rect 5356 13574 5358 13626
rect 5112 13572 5118 13574
rect 5174 13572 5198 13574
rect 5254 13572 5278 13574
rect 5334 13572 5358 13574
rect 5414 13572 5420 13574
rect 5112 13563 5420 13572
rect 5080 13524 5132 13530
rect 5000 13484 5080 13512
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 2780 12922 2832 12928
rect 3068 12940 3188 12968
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 10606 1808 12718
rect 2412 12436 2464 12442
rect 2516 12424 2544 12786
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2464 12396 2544 12424
rect 2412 12378 2464 12384
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11694 2544 12242
rect 2608 11694 2636 12718
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12102 2728 12582
rect 2792 12374 2820 12922
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2884 12442 2912 12718
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 3068 12238 3096 12940
rect 3988 12714 4016 13126
rect 4448 12986 4476 13194
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4724 12850 4752 13262
rect 4712 12844 4764 12850
rect 4764 12804 4844 12832
rect 4712 12786 4764 12792
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 12306 3188 12582
rect 3240 12368 3292 12374
rect 3240 12310 3292 12316
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2755 11996 3063 12005
rect 2755 11994 2761 11996
rect 2817 11994 2841 11996
rect 2897 11994 2921 11996
rect 2977 11994 3001 11996
rect 3057 11994 3063 11996
rect 2817 11942 2819 11994
rect 2999 11942 3001 11994
rect 2755 11940 2761 11942
rect 2817 11940 2841 11942
rect 2897 11940 2921 11942
rect 2977 11940 3001 11942
rect 3057 11940 3063 11942
rect 2755 11931 3063 11940
rect 3160 11898 3188 12038
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2976 11218 3004 11698
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 3068 11218 3096 11562
rect 3160 11354 3188 11834
rect 3252 11762 3280 12310
rect 4632 12306 4660 12650
rect 4816 12306 4844 12804
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3344 11558 3372 12174
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3988 11626 4016 12038
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1872 10538 1900 10950
rect 2755 10908 3063 10917
rect 2755 10906 2761 10908
rect 2817 10906 2841 10908
rect 2897 10906 2921 10908
rect 2977 10906 3001 10908
rect 3057 10906 3063 10908
rect 2817 10854 2819 10906
rect 2999 10854 3001 10906
rect 2755 10852 2761 10854
rect 2817 10852 2841 10854
rect 2897 10852 2921 10854
rect 2977 10852 3001 10854
rect 3057 10852 3063 10854
rect 2755 10843 3063 10852
rect 3160 10810 3188 11018
rect 3344 11014 3372 11494
rect 4080 11354 4108 12038
rect 4264 11354 4292 12242
rect 4908 12238 4936 12582
rect 5000 12442 5028 13484
rect 5080 13466 5132 13472
rect 5460 13394 5488 13670
rect 5448 13388 5500 13394
rect 5448 13330 5500 13336
rect 5460 12782 5488 13330
rect 5644 12986 5672 13874
rect 6932 13394 6960 13874
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5112 12540 5420 12549
rect 5112 12538 5118 12540
rect 5174 12538 5198 12540
rect 5254 12538 5278 12540
rect 5334 12538 5358 12540
rect 5414 12538 5420 12540
rect 5174 12486 5176 12538
rect 5356 12486 5358 12538
rect 5112 12484 5118 12486
rect 5174 12484 5198 12486
rect 5254 12484 5278 12486
rect 5334 12484 5358 12486
rect 5414 12484 5420 12486
rect 5112 12475 5420 12484
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4724 11830 4752 12174
rect 4908 11898 4936 12174
rect 5460 12102 5488 12582
rect 5644 12374 5672 12922
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4712 11824 4764 11830
rect 4712 11766 4764 11772
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4724 11268 4752 11766
rect 4804 11280 4856 11286
rect 4724 11240 4804 11268
rect 4804 11222 4856 11228
rect 4908 11014 4936 11834
rect 5644 11762 5672 12310
rect 6104 12238 6132 13126
rect 6920 12776 6972 12782
rect 6918 12744 6920 12753
rect 6972 12744 6974 12753
rect 6918 12679 6974 12688
rect 6092 12232 6144 12238
rect 6092 12174 6144 12180
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5828 11642 5856 11698
rect 6104 11694 6132 12174
rect 6092 11688 6144 11694
rect 5828 11614 6040 11642
rect 6092 11630 6144 11636
rect 6012 11558 6040 11614
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5112 11452 5420 11461
rect 5112 11450 5118 11452
rect 5174 11450 5198 11452
rect 5254 11450 5278 11452
rect 5334 11450 5358 11452
rect 5414 11450 5420 11452
rect 5174 11398 5176 11450
rect 5356 11398 5358 11450
rect 5112 11396 5118 11398
rect 5174 11396 5198 11398
rect 5254 11396 5278 11398
rect 5334 11396 5358 11398
rect 5414 11396 5420 11398
rect 5112 11387 5420 11396
rect 5460 11218 5488 11494
rect 6104 11354 6132 11630
rect 6644 11620 6696 11626
rect 6644 11562 6696 11568
rect 6656 11354 6684 11562
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 1860 10532 1912 10538
rect 1860 10474 1912 10480
rect 5112 10364 5420 10373
rect 5112 10362 5118 10364
rect 5174 10362 5198 10364
rect 5254 10362 5278 10364
rect 5334 10362 5358 10364
rect 5414 10362 5420 10364
rect 5174 10310 5176 10362
rect 5356 10310 5358 10362
rect 5112 10308 5118 10310
rect 5174 10308 5198 10310
rect 5254 10308 5278 10310
rect 5334 10308 5358 10310
rect 5414 10308 5420 10310
rect 5112 10299 5420 10308
rect 7024 10130 7052 18226
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7470 17436 7778 17445
rect 7470 17434 7476 17436
rect 7532 17434 7556 17436
rect 7612 17434 7636 17436
rect 7692 17434 7716 17436
rect 7772 17434 7778 17436
rect 7532 17382 7534 17434
rect 7714 17382 7716 17434
rect 7470 17380 7476 17382
rect 7532 17380 7556 17382
rect 7612 17380 7636 17382
rect 7692 17380 7716 17382
rect 7772 17380 7778 17382
rect 7470 17371 7778 17380
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7104 16516 7156 16522
rect 7104 16458 7156 16464
rect 7116 16114 7144 16458
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 7116 14482 7144 16050
rect 7208 15570 7236 17002
rect 7852 16794 7880 17002
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7944 16658 7972 17546
rect 8220 17134 8248 18226
rect 8312 18154 8340 18226
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8404 17882 8432 18022
rect 8392 17876 8444 17882
rect 8392 17818 8444 17824
rect 8392 17740 8444 17746
rect 8392 17682 8444 17688
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8312 16658 8340 17614
rect 8404 17542 8432 17682
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8404 16658 8432 17478
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 7470 16348 7778 16357
rect 7470 16346 7476 16348
rect 7532 16346 7556 16348
rect 7612 16346 7636 16348
rect 7692 16346 7716 16348
rect 7772 16346 7778 16348
rect 7532 16294 7534 16346
rect 7714 16294 7716 16346
rect 7470 16292 7476 16294
rect 7532 16292 7556 16294
rect 7612 16292 7636 16294
rect 7692 16292 7716 16294
rect 7772 16292 7778 16294
rect 7470 16283 7778 16292
rect 7840 15904 7892 15910
rect 7840 15846 7892 15852
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 14482 7236 15506
rect 7470 15260 7778 15269
rect 7470 15258 7476 15260
rect 7532 15258 7556 15260
rect 7612 15258 7636 15260
rect 7692 15258 7716 15260
rect 7772 15258 7778 15260
rect 7532 15206 7534 15258
rect 7714 15206 7716 15258
rect 7470 15204 7476 15206
rect 7532 15204 7556 15206
rect 7612 15204 7636 15206
rect 7692 15204 7716 15206
rect 7772 15204 7778 15206
rect 7470 15195 7778 15204
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7300 14482 7328 14758
rect 7852 14618 7880 15846
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7288 14476 7340 14482
rect 7288 14418 7340 14424
rect 7300 14006 7328 14418
rect 7470 14172 7778 14181
rect 7470 14170 7476 14172
rect 7532 14170 7556 14172
rect 7612 14170 7636 14172
rect 7692 14170 7716 14172
rect 7772 14170 7778 14172
rect 7532 14118 7534 14170
rect 7714 14118 7716 14170
rect 7470 14116 7476 14118
rect 7532 14116 7556 14118
rect 7612 14116 7636 14118
rect 7692 14116 7716 14118
rect 7772 14116 7778 14118
rect 7470 14107 7778 14116
rect 7288 14000 7340 14006
rect 7288 13942 7340 13948
rect 7944 13852 7972 16594
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8036 14362 8064 15982
rect 8036 14334 8248 14362
rect 7944 13824 8064 13852
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7470 13084 7778 13093
rect 7470 13082 7476 13084
rect 7532 13082 7556 13084
rect 7612 13082 7636 13084
rect 7692 13082 7716 13084
rect 7772 13082 7778 13084
rect 7532 13030 7534 13082
rect 7714 13030 7716 13082
rect 7470 13028 7476 13030
rect 7532 13028 7556 13030
rect 7612 13028 7636 13030
rect 7692 13028 7716 13030
rect 7772 13028 7778 13030
rect 7470 13019 7778 13028
rect 7852 12782 7880 13398
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7840 12776 7892 12782
rect 8036 12730 8064 13824
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7840 12718 7892 12724
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7116 12306 7144 12582
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7208 12102 7236 12718
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7470 11996 7778 12005
rect 7470 11994 7476 11996
rect 7532 11994 7556 11996
rect 7612 11994 7636 11996
rect 7692 11994 7716 11996
rect 7772 11994 7778 11996
rect 7532 11942 7534 11994
rect 7714 11942 7716 11994
rect 7470 11940 7476 11942
rect 7532 11940 7556 11942
rect 7612 11940 7636 11942
rect 7692 11940 7716 11942
rect 7772 11940 7778 11942
rect 7470 11931 7778 11940
rect 7852 11898 7880 12718
rect 7944 12702 8064 12730
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 7470 10908 7778 10917
rect 7470 10906 7476 10908
rect 7532 10906 7556 10908
rect 7612 10906 7636 10908
rect 7692 10906 7716 10908
rect 7772 10906 7778 10908
rect 7532 10854 7534 10906
rect 7714 10854 7716 10906
rect 7470 10852 7476 10854
rect 7532 10852 7556 10854
rect 7612 10852 7636 10854
rect 7692 10852 7716 10854
rect 7772 10852 7778 10854
rect 7470 10843 7778 10852
rect 7944 10606 7972 12702
rect 8128 12628 8156 12854
rect 8036 12600 8156 12628
rect 8036 10674 8064 12600
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7392 10130 7420 10542
rect 8220 10130 8248 14334
rect 8404 14278 8432 16594
rect 8496 16250 8524 17478
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 14618 8524 15846
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8404 13870 8432 14214
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8312 12986 8340 13262
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8404 12782 8432 13806
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8312 11286 8340 11630
rect 8404 11354 8432 11698
rect 8496 11354 8524 12174
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8300 11280 8352 11286
rect 8300 11222 8352 11228
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7380 10124 7432 10130
rect 7380 10066 7432 10072
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 2755 9820 3063 9829
rect 2755 9818 2761 9820
rect 2817 9818 2841 9820
rect 2897 9818 2921 9820
rect 2977 9818 3001 9820
rect 3057 9818 3063 9820
rect 2817 9766 2819 9818
rect 2999 9766 3001 9818
rect 2755 9764 2761 9766
rect 2817 9764 2841 9766
rect 2897 9764 2921 9766
rect 2977 9764 3001 9766
rect 3057 9764 3063 9766
rect 2755 9755 3063 9764
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5112 9276 5420 9285
rect 5112 9274 5118 9276
rect 5174 9274 5198 9276
rect 5254 9274 5278 9276
rect 5334 9274 5358 9276
rect 5414 9274 5420 9276
rect 5174 9222 5176 9274
rect 5356 9222 5358 9274
rect 5112 9220 5118 9222
rect 5174 9220 5198 9222
rect 5254 9220 5278 9222
rect 5334 9220 5358 9222
rect 5414 9220 5420 9222
rect 5112 9211 5420 9220
rect 2755 8732 3063 8741
rect 2755 8730 2761 8732
rect 2817 8730 2841 8732
rect 2897 8730 2921 8732
rect 2977 8730 3001 8732
rect 3057 8730 3063 8732
rect 2817 8678 2819 8730
rect 2999 8678 3001 8730
rect 2755 8676 2761 8678
rect 2817 8676 2841 8678
rect 2897 8676 2921 8678
rect 2977 8676 3001 8678
rect 3057 8676 3063 8678
rect 2755 8667 3063 8676
rect 5112 8188 5420 8197
rect 5112 8186 5118 8188
rect 5174 8186 5198 8188
rect 5254 8186 5278 8188
rect 5334 8186 5358 8188
rect 5414 8186 5420 8188
rect 5174 8134 5176 8186
rect 5356 8134 5358 8186
rect 5112 8132 5118 8134
rect 5174 8132 5198 8134
rect 5254 8132 5278 8134
rect 5334 8132 5358 8134
rect 5414 8132 5420 8134
rect 5112 8123 5420 8132
rect 2755 7644 3063 7653
rect 2755 7642 2761 7644
rect 2817 7642 2841 7644
rect 2897 7642 2921 7644
rect 2977 7642 3001 7644
rect 3057 7642 3063 7644
rect 2817 7590 2819 7642
rect 2999 7590 3001 7642
rect 2755 7588 2761 7590
rect 2817 7588 2841 7590
rect 2897 7588 2921 7590
rect 2977 7588 3001 7590
rect 3057 7588 3063 7590
rect 2755 7579 3063 7588
rect 5112 7100 5420 7109
rect 5112 7098 5118 7100
rect 5174 7098 5198 7100
rect 5254 7098 5278 7100
rect 5334 7098 5358 7100
rect 5414 7098 5420 7100
rect 5174 7046 5176 7098
rect 5356 7046 5358 7098
rect 5112 7044 5118 7046
rect 5174 7044 5198 7046
rect 5254 7044 5278 7046
rect 5334 7044 5358 7046
rect 5414 7044 5420 7046
rect 5112 7035 5420 7044
rect 2755 6556 3063 6565
rect 2755 6554 2761 6556
rect 2817 6554 2841 6556
rect 2897 6554 2921 6556
rect 2977 6554 3001 6556
rect 3057 6554 3063 6556
rect 2817 6502 2819 6554
rect 2999 6502 3001 6554
rect 2755 6500 2761 6502
rect 2817 6500 2841 6502
rect 2897 6500 2921 6502
rect 2977 6500 3001 6502
rect 3057 6500 3063 6502
rect 2755 6491 3063 6500
rect 5112 6012 5420 6021
rect 5112 6010 5118 6012
rect 5174 6010 5198 6012
rect 5254 6010 5278 6012
rect 5334 6010 5358 6012
rect 5414 6010 5420 6012
rect 5174 5958 5176 6010
rect 5356 5958 5358 6010
rect 5112 5956 5118 5958
rect 5174 5956 5198 5958
rect 5254 5956 5278 5958
rect 5334 5956 5358 5958
rect 5414 5956 5420 5958
rect 5112 5947 5420 5956
rect 2755 5468 3063 5477
rect 2755 5466 2761 5468
rect 2817 5466 2841 5468
rect 2897 5466 2921 5468
rect 2977 5466 3001 5468
rect 3057 5466 3063 5468
rect 2817 5414 2819 5466
rect 2999 5414 3001 5466
rect 2755 5412 2761 5414
rect 2817 5412 2841 5414
rect 2897 5412 2921 5414
rect 2977 5412 3001 5414
rect 3057 5412 3063 5414
rect 2755 5403 3063 5412
rect 5112 4924 5420 4933
rect 5112 4922 5118 4924
rect 5174 4922 5198 4924
rect 5254 4922 5278 4924
rect 5334 4922 5358 4924
rect 5414 4922 5420 4924
rect 5174 4870 5176 4922
rect 5356 4870 5358 4922
rect 5112 4868 5118 4870
rect 5174 4868 5198 4870
rect 5254 4868 5278 4870
rect 5334 4868 5358 4870
rect 5414 4868 5420 4870
rect 5112 4859 5420 4868
rect 2755 4380 3063 4389
rect 2755 4378 2761 4380
rect 2817 4378 2841 4380
rect 2897 4378 2921 4380
rect 2977 4378 3001 4380
rect 3057 4378 3063 4380
rect 2817 4326 2819 4378
rect 2999 4326 3001 4378
rect 2755 4324 2761 4326
rect 2817 4324 2841 4326
rect 2897 4324 2921 4326
rect 2977 4324 3001 4326
rect 3057 4324 3063 4326
rect 2755 4315 3063 4324
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 1216 3528 1268 3534
rect 1216 3470 1268 3476
rect 1228 400 1256 3470
rect 2755 3292 3063 3301
rect 2755 3290 2761 3292
rect 2817 3290 2841 3292
rect 2897 3290 2921 3292
rect 2977 3290 3001 3292
rect 3057 3290 3063 3292
rect 2817 3238 2819 3290
rect 2999 3238 3001 3290
rect 2755 3236 2761 3238
rect 2817 3236 2841 3238
rect 2897 3236 2921 3238
rect 2977 3236 3001 3238
rect 3057 3236 3063 3238
rect 2755 3227 3063 3236
rect 2755 2204 3063 2213
rect 2755 2202 2761 2204
rect 2817 2202 2841 2204
rect 2897 2202 2921 2204
rect 2977 2202 3001 2204
rect 3057 2202 3063 2204
rect 2817 2150 2819 2202
rect 2999 2150 3001 2202
rect 2755 2148 2761 2150
rect 2817 2148 2841 2150
rect 2897 2148 2921 2150
rect 2977 2148 3001 2150
rect 3057 2148 3063 2150
rect 2755 2139 3063 2148
rect 2755 1116 3063 1125
rect 2755 1114 2761 1116
rect 2817 1114 2841 1116
rect 2897 1114 2921 1116
rect 2977 1114 3001 1116
rect 3057 1114 3063 1116
rect 2817 1062 2819 1114
rect 2999 1062 3001 1114
rect 2755 1060 2761 1062
rect 2817 1060 2841 1062
rect 2897 1060 2921 1062
rect 2977 1060 3001 1062
rect 3057 1060 3063 1062
rect 2755 1051 3063 1060
rect 3712 400 3740 4082
rect 5112 3836 5420 3845
rect 5112 3834 5118 3836
rect 5174 3834 5198 3836
rect 5254 3834 5278 3836
rect 5334 3834 5358 3836
rect 5414 3834 5420 3836
rect 5174 3782 5176 3834
rect 5356 3782 5358 3834
rect 5112 3780 5118 3782
rect 5174 3780 5198 3782
rect 5254 3780 5278 3782
rect 5334 3780 5358 3782
rect 5414 3780 5420 3782
rect 5112 3771 5420 3780
rect 5112 2748 5420 2757
rect 5112 2746 5118 2748
rect 5174 2746 5198 2748
rect 5254 2746 5278 2748
rect 5334 2746 5358 2748
rect 5414 2746 5420 2748
rect 5174 2694 5176 2746
rect 5356 2694 5358 2746
rect 5112 2692 5118 2694
rect 5174 2692 5198 2694
rect 5254 2692 5278 2694
rect 5334 2692 5358 2694
rect 5414 2692 5420 2694
rect 5112 2683 5420 2692
rect 5112 1660 5420 1669
rect 5112 1658 5118 1660
rect 5174 1658 5198 1660
rect 5254 1658 5278 1660
rect 5334 1658 5358 1660
rect 5414 1658 5420 1660
rect 5174 1606 5176 1658
rect 5356 1606 5358 1658
rect 5112 1604 5118 1606
rect 5174 1604 5198 1606
rect 5254 1604 5278 1606
rect 5334 1604 5358 1606
rect 5414 1604 5420 1606
rect 5112 1595 5420 1604
rect 5112 572 5420 581
rect 5112 570 5118 572
rect 5174 570 5198 572
rect 5254 570 5278 572
rect 5334 570 5358 572
rect 5414 570 5420 572
rect 5174 518 5176 570
rect 5356 518 5358 570
rect 5112 516 5118 518
rect 5174 516 5198 518
rect 5254 516 5278 518
rect 5334 516 5358 518
rect 5414 516 5420 518
rect 5112 507 5420 516
rect 6196 400 6224 9318
rect 7392 9178 7420 9862
rect 7470 9820 7778 9829
rect 7470 9818 7476 9820
rect 7532 9818 7556 9820
rect 7612 9818 7636 9820
rect 7692 9818 7716 9820
rect 7772 9818 7778 9820
rect 7532 9766 7534 9818
rect 7714 9766 7716 9818
rect 7470 9764 7476 9766
rect 7532 9764 7556 9766
rect 7612 9764 7636 9766
rect 7692 9764 7716 9766
rect 7772 9764 7778 9766
rect 7470 9755 7778 9764
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7472 9376 7524 9382
rect 7472 9318 7524 9324
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7484 9042 7512 9318
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 7668 8906 7696 9386
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7470 8732 7778 8741
rect 7470 8730 7476 8732
rect 7532 8730 7556 8732
rect 7612 8730 7636 8732
rect 7692 8730 7716 8732
rect 7772 8730 7778 8732
rect 7532 8678 7534 8730
rect 7714 8678 7716 8730
rect 7470 8676 7476 8678
rect 7532 8676 7556 8678
rect 7612 8676 7636 8678
rect 7692 8676 7716 8678
rect 7772 8676 7778 8678
rect 7470 8667 7778 8676
rect 7470 7644 7778 7653
rect 7470 7642 7476 7644
rect 7532 7642 7556 7644
rect 7612 7642 7636 7644
rect 7692 7642 7716 7644
rect 7772 7642 7778 7644
rect 7532 7590 7534 7642
rect 7714 7590 7716 7642
rect 7470 7588 7476 7590
rect 7532 7588 7556 7590
rect 7612 7588 7636 7590
rect 7692 7588 7716 7590
rect 7772 7588 7778 7590
rect 7470 7579 7778 7588
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6564 3534 6592 7210
rect 8312 7206 8340 10406
rect 8404 9586 8432 10542
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8404 8430 8432 9522
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 7478 8432 8366
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7470 6556 7778 6565
rect 7470 6554 7476 6556
rect 7532 6554 7556 6556
rect 7612 6554 7636 6556
rect 7692 6554 7716 6556
rect 7772 6554 7778 6556
rect 7532 6502 7534 6554
rect 7714 6502 7716 6554
rect 7470 6500 7476 6502
rect 7532 6500 7556 6502
rect 7612 6500 7636 6502
rect 7692 6500 7716 6502
rect 7772 6500 7778 6502
rect 7470 6491 7778 6500
rect 8404 6254 8432 7414
rect 8496 7342 8524 7686
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8588 6866 8616 18566
rect 8680 15688 8708 18906
rect 9140 18902 9168 19600
rect 9827 19068 10135 19077
rect 9827 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10073 19068
rect 10129 19066 10135 19068
rect 9889 19014 9891 19066
rect 10071 19014 10073 19066
rect 9827 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10073 19014
rect 10129 19012 10135 19014
rect 9827 19003 10135 19012
rect 9128 18896 9180 18902
rect 9128 18838 9180 18844
rect 10796 18834 10824 19600
rect 12452 18834 12480 19600
rect 14108 18834 14136 19600
rect 14542 19068 14850 19077
rect 14542 19066 14548 19068
rect 14604 19066 14628 19068
rect 14684 19066 14708 19068
rect 14764 19066 14788 19068
rect 14844 19066 14850 19068
rect 14604 19014 14606 19066
rect 14786 19014 14788 19066
rect 14542 19012 14548 19014
rect 14604 19012 14628 19014
rect 14684 19012 14708 19014
rect 14764 19012 14788 19014
rect 14844 19012 14850 19014
rect 14542 19003 14850 19012
rect 15764 18834 15792 19600
rect 17420 18834 17448 19600
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 14096 18828 14148 18834
rect 14096 18770 14148 18776
rect 15752 18828 15804 18834
rect 15752 18770 15804 18776
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9220 18692 9272 18698
rect 9220 18634 9272 18640
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 18154 8984 18226
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 9048 17882 9076 18294
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8760 16720 8812 16726
rect 8864 16697 8892 17274
rect 8760 16662 8812 16668
rect 8850 16688 8906 16697
rect 8772 16114 8800 16662
rect 8850 16623 8906 16632
rect 8864 16454 8892 16623
rect 9140 16522 9168 18022
rect 9232 16658 9260 18634
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9324 17542 9352 18362
rect 9404 18216 9456 18222
rect 9508 18170 9536 18566
rect 9600 18222 9628 18702
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9456 18164 9536 18170
rect 9404 18158 9536 18164
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9416 18142 9536 18158
rect 9508 17746 9536 18142
rect 9692 17746 9720 18634
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 9827 17980 10135 17989
rect 9827 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10073 17980
rect 10129 17978 10135 17980
rect 9889 17926 9891 17978
rect 10071 17926 10073 17978
rect 9827 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10073 17926
rect 10129 17924 10135 17926
rect 9827 17915 10135 17924
rect 10612 17746 10640 18566
rect 12185 18524 12493 18533
rect 12185 18522 12191 18524
rect 12247 18522 12271 18524
rect 12327 18522 12351 18524
rect 12407 18522 12431 18524
rect 12487 18522 12493 18524
rect 12247 18470 12249 18522
rect 12429 18470 12431 18522
rect 12185 18468 12191 18470
rect 12247 18468 12271 18470
rect 12327 18468 12351 18470
rect 12407 18468 12431 18470
rect 12487 18468 12493 18470
rect 12185 18459 12493 18468
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8760 16108 8812 16114
rect 8760 16050 8812 16056
rect 8956 16046 8984 16390
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 9036 16040 9088 16046
rect 9036 15982 9088 15988
rect 8680 15660 8800 15688
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8680 15473 8708 15506
rect 8666 15464 8722 15473
rect 8666 15399 8722 15408
rect 8772 14346 8800 15660
rect 9048 15162 9076 15982
rect 9232 15570 9260 16186
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9416 15638 9444 16118
rect 9404 15632 9456 15638
rect 9404 15574 9456 15580
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14618 8984 14826
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 9048 13462 9076 15098
rect 9140 14958 9168 15438
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8680 11218 8708 12854
rect 9048 12850 9076 13398
rect 9140 13394 9168 14894
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9416 12782 9444 13398
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 8956 12646 8984 12718
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 8852 11620 8904 11626
rect 8852 11562 8904 11568
rect 8864 11218 8892 11562
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8956 9110 8984 12582
rect 9416 12306 9444 12582
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9508 12186 9536 17478
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9692 16794 9720 17002
rect 9827 16892 10135 16901
rect 9827 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10073 16892
rect 10129 16890 10135 16892
rect 9889 16838 9891 16890
rect 10071 16838 10073 16890
rect 9827 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10073 16838
rect 10129 16836 10135 16838
rect 9827 16827 10135 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9956 16720 10008 16726
rect 9954 16688 9956 16697
rect 10008 16688 10010 16697
rect 10244 16658 10272 17682
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 17542 11468 17614
rect 10416 17536 10468 17542
rect 10416 17478 10468 17484
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 9954 16623 10010 16632
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9600 16046 9628 16458
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9692 12986 9720 16526
rect 10428 15978 10456 17478
rect 11440 16726 11468 17478
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10888 16250 10916 16390
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 9827 15804 10135 15813
rect 9827 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10073 15804
rect 10129 15802 10135 15804
rect 9889 15750 9891 15802
rect 10071 15750 10073 15802
rect 9827 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10073 15750
rect 10129 15748 10135 15750
rect 9827 15739 10135 15748
rect 10428 15586 10456 15914
rect 10520 15706 10548 16186
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10428 15558 10548 15586
rect 9827 14716 10135 14725
rect 9827 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10073 14716
rect 10129 14714 10135 14716
rect 9889 14662 9891 14714
rect 10071 14662 10073 14714
rect 9827 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10073 14662
rect 10129 14660 10135 14662
rect 9827 14651 10135 14660
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 9827 13628 10135 13637
rect 9827 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10073 13628
rect 10129 13626 10135 13628
rect 9889 13574 9891 13626
rect 10071 13574 10073 13626
rect 9827 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10073 13574
rect 10129 13572 10135 13574
rect 9827 13563 10135 13572
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12986 9996 13330
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10244 12782 10272 13670
rect 9680 12776 9732 12782
rect 9586 12744 9642 12753
rect 9680 12718 9732 12724
rect 10232 12776 10284 12782
rect 10232 12718 10284 12724
rect 10324 12776 10376 12782
rect 10324 12718 10376 12724
rect 9586 12679 9642 12688
rect 9416 12158 9536 12186
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10606 9076 10950
rect 9036 10600 9088 10606
rect 9036 10542 9088 10548
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8392 6248 8444 6254
rect 8392 6190 8444 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 7470 5468 7778 5477
rect 7470 5466 7476 5468
rect 7532 5466 7556 5468
rect 7612 5466 7636 5468
rect 7692 5466 7716 5468
rect 7772 5466 7778 5468
rect 7532 5414 7534 5466
rect 7714 5414 7716 5466
rect 7470 5412 7476 5414
rect 7532 5412 7556 5414
rect 7612 5412 7636 5414
rect 7692 5412 7716 5414
rect 7772 5412 7778 5414
rect 7470 5403 7778 5412
rect 7470 4380 7778 4389
rect 7470 4378 7476 4380
rect 7532 4378 7556 4380
rect 7612 4378 7636 4380
rect 7692 4378 7716 4380
rect 7772 4378 7778 4380
rect 7532 4326 7534 4378
rect 7714 4326 7716 4378
rect 7470 4324 7476 4326
rect 7532 4324 7556 4326
rect 7612 4324 7636 4326
rect 7692 4324 7716 4326
rect 7772 4324 7778 4326
rect 7470 4315 7778 4324
rect 8496 4146 8524 6054
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 7470 3292 7778 3301
rect 7470 3290 7476 3292
rect 7532 3290 7556 3292
rect 7612 3290 7636 3292
rect 7692 3290 7716 3292
rect 7772 3290 7778 3292
rect 7532 3238 7534 3290
rect 7714 3238 7716 3290
rect 7470 3236 7476 3238
rect 7532 3236 7556 3238
rect 7612 3236 7636 3238
rect 7692 3236 7716 3238
rect 7772 3236 7778 3238
rect 7470 3227 7778 3236
rect 7470 2204 7778 2213
rect 7470 2202 7476 2204
rect 7532 2202 7556 2204
rect 7612 2202 7636 2204
rect 7692 2202 7716 2204
rect 7772 2202 7778 2204
rect 7532 2150 7534 2202
rect 7714 2150 7716 2202
rect 7470 2148 7476 2150
rect 7532 2148 7556 2150
rect 7612 2148 7636 2150
rect 7692 2148 7716 2150
rect 7772 2148 7778 2150
rect 7470 2139 7778 2148
rect 7470 1116 7778 1125
rect 7470 1114 7476 1116
rect 7532 1114 7556 1116
rect 7612 1114 7636 1116
rect 7692 1114 7716 1116
rect 7772 1114 7778 1116
rect 7532 1062 7534 1114
rect 7714 1062 7716 1114
rect 7470 1060 7476 1062
rect 7532 1060 7556 1062
rect 7612 1060 7636 1062
rect 7692 1060 7716 1062
rect 7772 1060 7778 1062
rect 7470 1051 7778 1060
rect 8680 400 8708 8502
rect 8864 8362 8892 8774
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8956 7342 8984 9046
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8956 6934 8984 7278
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8956 6458 8984 6870
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5778 9352 6190
rect 9416 6118 9444 12158
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11286 9536 12038
rect 9600 11558 9628 12679
rect 9692 12434 9720 12718
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9827 12540 10135 12549
rect 9827 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10073 12540
rect 10129 12538 10135 12540
rect 9889 12486 9891 12538
rect 10071 12486 10073 12538
rect 9827 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10073 12486
rect 10129 12484 10135 12486
rect 9827 12475 10135 12484
rect 9692 12406 9904 12434
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11694 9812 12174
rect 9876 12170 9904 12406
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9588 11552 9640 11558
rect 9784 11540 9812 11630
rect 9876 11626 9904 12106
rect 10152 11762 10180 12310
rect 10244 12238 10272 12582
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9588 11494 9640 11500
rect 9692 11512 9812 11540
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9508 10810 9536 11086
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9508 10130 9536 10746
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9382 9536 9862
rect 9600 9602 9628 11494
rect 9692 11218 9720 11512
rect 9827 11452 10135 11461
rect 9827 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10073 11452
rect 10129 11450 10135 11452
rect 9889 11398 9891 11450
rect 10071 11398 10073 11450
rect 9827 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10073 11398
rect 10129 11396 10135 11398
rect 9827 11387 10135 11396
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 9784 11218 9812 11290
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9692 10742 9720 11154
rect 10244 11098 10272 11290
rect 10336 11218 10364 12718
rect 10520 12594 10548 15558
rect 10612 15366 10640 15982
rect 11164 15570 11192 16594
rect 11256 16046 11284 16594
rect 11244 16040 11296 16046
rect 11244 15982 11296 15988
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15706 11376 15982
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10612 14890 10640 15302
rect 10600 14884 10652 14890
rect 10600 14826 10652 14832
rect 10428 12566 10548 12594
rect 10428 11558 10456 12566
rect 10612 12434 10640 14826
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10520 12406 10640 12434
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10416 11280 10468 11286
rect 10520 11268 10548 12406
rect 10598 11792 10654 11801
rect 10598 11727 10654 11736
rect 10612 11694 10640 11727
rect 10704 11694 10732 12854
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10468 11240 10548 11268
rect 10416 11222 10468 11228
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10152 11082 10272 11098
rect 10140 11076 10272 11082
rect 10192 11070 10272 11076
rect 10140 11018 10192 11024
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9827 10364 10135 10373
rect 9827 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10073 10364
rect 10129 10362 10135 10364
rect 9889 10310 9891 10362
rect 10071 10310 10073 10362
rect 9827 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10073 10310
rect 10129 10308 10135 10310
rect 9827 10299 10135 10308
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9600 9574 9720 9602
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9508 9042 9536 9318
rect 9692 9058 9720 9574
rect 9784 9518 9812 9998
rect 9968 9722 9996 10066
rect 10152 9994 10180 10066
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9968 9518 9996 9658
rect 10046 9616 10102 9625
rect 10046 9551 10102 9560
rect 10060 9518 10088 9551
rect 10152 9518 10180 9930
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 9827 9276 10135 9285
rect 9827 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10073 9276
rect 10129 9274 10135 9276
rect 9889 9222 9891 9274
rect 10071 9222 10073 9274
rect 9827 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10073 9222
rect 10129 9220 10135 9222
rect 9827 9211 10135 9220
rect 9496 9036 9548 9042
rect 9692 9030 9812 9058
rect 10244 9042 10272 9658
rect 9496 8978 9548 8984
rect 9508 8022 9536 8978
rect 9784 8362 9812 9030
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 10336 8838 10364 9998
rect 10428 9382 10456 11222
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10416 8968 10468 8974
rect 10612 8956 10640 11494
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10468 8928 10640 8956
rect 10416 8910 10468 8916
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9827 8188 10135 8197
rect 9827 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10073 8188
rect 10129 8186 10135 8188
rect 9889 8134 9891 8186
rect 10071 8134 10073 8186
rect 9827 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10073 8134
rect 10129 8132 10135 8134
rect 9827 8123 10135 8132
rect 10336 8090 10364 8774
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9508 7342 9536 7958
rect 9876 7342 9904 8026
rect 9496 7336 9548 7342
rect 9864 7336 9916 7342
rect 9496 7278 9548 7284
rect 9692 7296 9864 7324
rect 9508 6934 9536 7278
rect 9692 7002 9720 7296
rect 9864 7278 9916 7284
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 9827 7100 10135 7109
rect 9827 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10073 7100
rect 10129 7098 10135 7100
rect 9889 7046 9891 7098
rect 10071 7046 10073 7098
rect 9827 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10073 7046
rect 10129 7044 10135 7046
rect 9827 7035 10135 7044
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9600 6186 9628 6598
rect 9968 6254 9996 6598
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9827 6012 10135 6021
rect 9827 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10073 6012
rect 10129 6010 10135 6012
rect 9889 5958 9891 6010
rect 10071 5958 10073 6010
rect 9827 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10073 5958
rect 10129 5956 10135 5958
rect 9827 5947 10135 5956
rect 10244 5794 10272 6326
rect 10336 6254 10364 7142
rect 10704 6254 10732 10202
rect 10796 9625 10824 14282
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 12782 10916 13670
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10980 12850 11008 13126
rect 11072 12986 11100 13738
rect 11164 13530 11192 15370
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11440 14550 11468 15302
rect 11532 15162 11560 16730
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 11624 16046 11652 16390
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11716 15570 11744 17682
rect 12185 17436 12493 17445
rect 12185 17434 12191 17436
rect 12247 17434 12271 17436
rect 12327 17434 12351 17436
rect 12407 17434 12431 17436
rect 12487 17434 12493 17436
rect 12247 17382 12249 17434
rect 12429 17382 12431 17434
rect 12185 17380 12191 17382
rect 12247 17380 12271 17382
rect 12327 17380 12351 17382
rect 12407 17380 12431 17382
rect 12487 17380 12493 17382
rect 12185 17371 12493 17380
rect 11808 16658 12112 16674
rect 11796 16652 12124 16658
rect 11848 16646 12072 16652
rect 11796 16594 11848 16600
rect 12072 16594 12124 16600
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 16454 12020 16526
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11808 15570 11836 16390
rect 11992 15570 12020 16390
rect 12185 16348 12493 16357
rect 12185 16346 12191 16348
rect 12247 16346 12271 16348
rect 12327 16346 12351 16348
rect 12407 16346 12431 16348
rect 12487 16346 12493 16348
rect 12247 16294 12249 16346
rect 12429 16294 12431 16346
rect 12185 16292 12191 16294
rect 12247 16292 12271 16294
rect 12327 16292 12351 16294
rect 12407 16292 12431 16294
rect 12487 16292 12493 16294
rect 12185 16283 12493 16292
rect 12544 16250 12572 18566
rect 14464 18080 14516 18086
rect 14464 18022 14516 18028
rect 14476 17814 14504 18022
rect 14542 17980 14850 17989
rect 14542 17978 14548 17980
rect 14604 17978 14628 17980
rect 14684 17978 14708 17980
rect 14764 17978 14788 17980
rect 14844 17978 14850 17980
rect 14604 17926 14606 17978
rect 14786 17926 14788 17978
rect 14542 17924 14548 17926
rect 14604 17924 14628 17926
rect 14684 17924 14708 17926
rect 14764 17924 14788 17926
rect 14844 17924 14850 17926
rect 14542 17915 14850 17924
rect 14464 17808 14516 17814
rect 14464 17750 14516 17756
rect 16132 17678 16160 18566
rect 16776 18222 16804 18566
rect 16900 18524 17208 18533
rect 16900 18522 16906 18524
rect 16962 18522 16986 18524
rect 17042 18522 17066 18524
rect 17122 18522 17146 18524
rect 17202 18522 17208 18524
rect 16962 18470 16964 18522
rect 17144 18470 17146 18522
rect 16900 18468 16906 18470
rect 16962 18468 16986 18470
rect 17042 18468 17066 18470
rect 17122 18468 17146 18470
rect 17202 18468 17208 18470
rect 16900 18459 17208 18468
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16684 17814 16712 18022
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12256 15904 12308 15910
rect 12256 15846 12308 15852
rect 12268 15570 12296 15846
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11520 15156 11572 15162
rect 11520 15098 11572 15104
rect 11900 14890 11928 15302
rect 12185 15260 12493 15269
rect 12185 15258 12191 15260
rect 12247 15258 12271 15260
rect 12327 15258 12351 15260
rect 12407 15258 12431 15260
rect 12487 15258 12493 15260
rect 12247 15206 12249 15258
rect 12429 15206 12431 15258
rect 12185 15204 12191 15206
rect 12247 15204 12271 15206
rect 12327 15204 12351 15206
rect 12407 15204 12431 15206
rect 12487 15204 12493 15206
rect 12185 15195 12493 15204
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 11624 14482 11652 14826
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11612 14476 11664 14482
rect 11532 14436 11612 14464
rect 11532 13802 11560 14436
rect 11612 14418 11664 14424
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11624 13376 11652 14214
rect 11716 14074 11744 14282
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11900 13870 11928 14350
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13394 11836 13670
rect 11992 13394 12020 14418
rect 12084 14074 12112 14486
rect 12544 14482 12572 15982
rect 12636 15570 12664 16526
rect 13556 16114 13584 17614
rect 16900 17436 17208 17445
rect 16900 17434 16906 17436
rect 16962 17434 16986 17436
rect 17042 17434 17066 17436
rect 17122 17434 17146 17436
rect 17202 17434 17208 17436
rect 16962 17382 16964 17434
rect 17144 17382 17146 17434
rect 16900 17380 16906 17382
rect 16962 17380 16986 17382
rect 17042 17380 17066 17382
rect 17122 17380 17146 17382
rect 17202 17380 17208 17382
rect 16900 17371 17208 17380
rect 14542 16892 14850 16901
rect 14542 16890 14548 16892
rect 14604 16890 14628 16892
rect 14684 16890 14708 16892
rect 14764 16890 14788 16892
rect 14844 16890 14850 16892
rect 14604 16838 14606 16890
rect 14786 16838 14788 16890
rect 14542 16836 14548 16838
rect 14604 16836 14628 16838
rect 14684 16836 14708 16838
rect 14764 16836 14788 16838
rect 14844 16836 14850 16838
rect 14542 16827 14850 16836
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15706 13860 15982
rect 15212 15910 15240 16526
rect 16900 16348 17208 16357
rect 16900 16346 16906 16348
rect 16962 16346 16986 16348
rect 17042 16346 17066 16348
rect 17122 16346 17146 16348
rect 17202 16346 17208 16348
rect 16962 16294 16964 16346
rect 17144 16294 17146 16346
rect 16900 16292 16906 16294
rect 16962 16292 16986 16294
rect 17042 16292 17066 16294
rect 17122 16292 17146 16294
rect 17202 16292 17208 16294
rect 16900 16283 17208 16292
rect 19076 16017 19104 19600
rect 19257 19068 19565 19077
rect 19257 19066 19263 19068
rect 19319 19066 19343 19068
rect 19399 19066 19423 19068
rect 19479 19066 19503 19068
rect 19559 19066 19565 19068
rect 19319 19014 19321 19066
rect 19501 19014 19503 19066
rect 19257 19012 19263 19014
rect 19319 19012 19343 19014
rect 19399 19012 19423 19014
rect 19479 19012 19503 19014
rect 19559 19012 19565 19014
rect 19257 19003 19565 19012
rect 19257 17980 19565 17989
rect 19257 17978 19263 17980
rect 19319 17978 19343 17980
rect 19399 17978 19423 17980
rect 19479 17978 19503 17980
rect 19559 17978 19565 17980
rect 19319 17926 19321 17978
rect 19501 17926 19503 17978
rect 19257 17924 19263 17926
rect 19319 17924 19343 17926
rect 19399 17924 19423 17926
rect 19479 17924 19503 17926
rect 19559 17924 19565 17926
rect 19257 17915 19565 17924
rect 19257 16892 19565 16901
rect 19257 16890 19263 16892
rect 19319 16890 19343 16892
rect 19399 16890 19423 16892
rect 19479 16890 19503 16892
rect 19559 16890 19565 16892
rect 19319 16838 19321 16890
rect 19501 16838 19503 16890
rect 19257 16836 19263 16838
rect 19319 16836 19343 16838
rect 19399 16836 19423 16838
rect 19479 16836 19503 16838
rect 19559 16836 19565 16838
rect 19257 16827 19565 16836
rect 19062 16008 19118 16017
rect 19062 15943 19118 15952
rect 14832 15904 14884 15910
rect 15200 15904 15252 15910
rect 14884 15864 14964 15892
rect 14832 15846 14884 15852
rect 14542 15804 14850 15813
rect 14542 15802 14548 15804
rect 14604 15802 14628 15804
rect 14684 15802 14708 15804
rect 14764 15802 14788 15804
rect 14844 15802 14850 15804
rect 14604 15750 14606 15802
rect 14786 15750 14788 15802
rect 14542 15748 14548 15750
rect 14604 15748 14628 15750
rect 14684 15748 14708 15750
rect 14764 15748 14788 15750
rect 14844 15748 14850 15750
rect 14542 15739 14850 15748
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12912 15162 12940 15506
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 14936 14958 14964 15864
rect 15200 15846 15252 15852
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14542 14716 14850 14725
rect 14542 14714 14548 14716
rect 14604 14714 14628 14716
rect 14684 14714 14708 14716
rect 14764 14714 14788 14716
rect 14844 14714 14850 14716
rect 14604 14662 14606 14714
rect 14786 14662 14788 14714
rect 14542 14660 14548 14662
rect 14604 14660 14628 14662
rect 14684 14660 14708 14662
rect 14764 14660 14788 14662
rect 14844 14660 14850 14662
rect 14542 14651 14850 14660
rect 14936 14482 14964 14894
rect 15212 14890 15240 15846
rect 19257 15804 19565 15813
rect 19257 15802 19263 15804
rect 19319 15802 19343 15804
rect 19399 15802 19423 15804
rect 19479 15802 19503 15804
rect 19559 15802 19565 15804
rect 19319 15750 19321 15802
rect 19501 15750 19503 15802
rect 19257 15748 19263 15750
rect 19319 15748 19343 15750
rect 19399 15748 19423 15750
rect 19479 15748 19503 15750
rect 19559 15748 19565 15750
rect 19257 15739 19565 15748
rect 16900 15260 17208 15269
rect 16900 15258 16906 15260
rect 16962 15258 16986 15260
rect 17042 15258 17066 15260
rect 17122 15258 17146 15260
rect 17202 15258 17208 15260
rect 16962 15206 16964 15258
rect 17144 15206 17146 15258
rect 16900 15204 16906 15206
rect 16962 15204 16986 15206
rect 17042 15204 17066 15206
rect 17122 15204 17146 15206
rect 17202 15204 17208 15206
rect 16900 15195 17208 15204
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 14924 14476 14976 14482
rect 15108 14476 15160 14482
rect 14924 14418 14976 14424
rect 15028 14436 15108 14464
rect 12185 14172 12493 14181
rect 12185 14170 12191 14172
rect 12247 14170 12271 14172
rect 12327 14170 12351 14172
rect 12407 14170 12431 14172
rect 12487 14170 12493 14172
rect 12247 14118 12249 14170
rect 12429 14118 12431 14170
rect 12185 14116 12191 14118
rect 12247 14116 12271 14118
rect 12327 14116 12351 14118
rect 12407 14116 12431 14118
rect 12487 14116 12493 14118
rect 12185 14107 12493 14116
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11704 13388 11756 13394
rect 11624 13348 11704 13376
rect 11704 13330 11756 13336
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12844 11020 12850
rect 10968 12786 11020 12792
rect 11348 12782 11376 13194
rect 11716 12918 11744 13330
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12084 12986 12112 13262
rect 12185 13084 12493 13093
rect 12185 13082 12191 13084
rect 12247 13082 12271 13084
rect 12327 13082 12351 13084
rect 12407 13082 12431 13084
rect 12487 13082 12493 13084
rect 12247 13030 12249 13082
rect 12429 13030 12431 13082
rect 12185 13028 12191 13030
rect 12247 13028 12271 13030
rect 12327 13028 12351 13030
rect 12407 13028 12431 13030
rect 12487 13028 12493 13030
rect 12185 13019 12493 13028
rect 12544 12986 12572 14418
rect 12728 14074 12756 14418
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12820 13870 12848 14214
rect 13832 13870 13860 14214
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 11704 12912 11756 12918
rect 11704 12854 11756 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11518 12744 11574 12753
rect 10888 12238 10916 12718
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10980 12442 11008 12650
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10888 11694 10916 12038
rect 11072 11898 11100 12242
rect 11060 11892 11112 11898
rect 11060 11834 11112 11840
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 11348 11218 11376 12718
rect 11518 12679 11520 12688
rect 11572 12679 11574 12688
rect 11520 12650 11572 12656
rect 12084 12374 12112 12922
rect 12636 12442 12664 13806
rect 14542 13628 14850 13637
rect 14542 13626 14548 13628
rect 14604 13626 14628 13628
rect 14684 13626 14708 13628
rect 14764 13626 14788 13628
rect 14844 13626 14850 13628
rect 14604 13574 14606 13626
rect 14786 13574 14788 13626
rect 14542 13572 14548 13574
rect 14604 13572 14628 13574
rect 14684 13572 14708 13574
rect 14764 13572 14788 13574
rect 14844 13572 14850 13574
rect 14542 13563 14850 13572
rect 15028 13530 15056 14436
rect 15108 14418 15160 14424
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13360 12708 13412 12714
rect 13360 12650 13412 12656
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 13372 12306 13400 12650
rect 13740 12306 13768 13126
rect 15028 12782 15056 13466
rect 15120 13394 15148 13806
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15120 12782 15148 13330
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 14542 12540 14850 12549
rect 14542 12538 14548 12540
rect 14604 12538 14628 12540
rect 14684 12538 14708 12540
rect 14764 12538 14788 12540
rect 14844 12538 14850 12540
rect 14604 12486 14606 12538
rect 14786 12486 14788 12538
rect 14542 12484 14548 12486
rect 14604 12484 14628 12486
rect 14684 12484 14708 12486
rect 14764 12484 14788 12486
rect 14844 12484 14850 12486
rect 14542 12475 14850 12484
rect 15028 12374 15056 12718
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 12185 11996 12493 12005
rect 12185 11994 12191 11996
rect 12247 11994 12271 11996
rect 12327 11994 12351 11996
rect 12407 11994 12431 11996
rect 12487 11994 12493 11996
rect 12247 11942 12249 11994
rect 12429 11942 12431 11994
rect 12185 11940 12191 11942
rect 12247 11940 12271 11942
rect 12327 11940 12351 11942
rect 12407 11940 12431 11942
rect 12487 11940 12493 11942
rect 12185 11931 12493 11940
rect 13372 11694 13400 12242
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 12636 11218 12664 11630
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10130 11284 10678
rect 11348 10674 11376 11154
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11440 10606 11468 11086
rect 12185 10908 12493 10917
rect 12185 10906 12191 10908
rect 12247 10906 12271 10908
rect 12327 10906 12351 10908
rect 12407 10906 12431 10908
rect 12487 10906 12493 10908
rect 12247 10854 12249 10906
rect 12429 10854 12431 10906
rect 12185 10852 12191 10854
rect 12247 10852 12271 10854
rect 12327 10852 12351 10854
rect 12407 10852 12431 10854
rect 12487 10852 12493 10854
rect 12185 10843 12493 10852
rect 12636 10606 12664 11154
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 11428 10600 11480 10606
rect 11428 10542 11480 10548
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 10782 9616 10838 9625
rect 10782 9551 10838 9560
rect 11256 9518 11284 10066
rect 11440 9586 11468 10542
rect 12636 10130 12664 10542
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12185 9820 12493 9829
rect 12185 9818 12191 9820
rect 12247 9818 12271 9820
rect 12327 9818 12351 9820
rect 12407 9818 12431 9820
rect 12487 9818 12493 9820
rect 12247 9766 12249 9818
rect 12429 9766 12431 9818
rect 12185 9764 12191 9766
rect 12247 9764 12271 9766
rect 12327 9764 12351 9766
rect 12407 9764 12431 9766
rect 12487 9764 12493 9766
rect 12185 9755 12493 9764
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11532 9042 11560 9114
rect 11900 9042 11928 9318
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 11532 7342 11560 8978
rect 11808 8634 11836 8978
rect 12185 8732 12493 8741
rect 12185 8730 12191 8732
rect 12247 8730 12271 8732
rect 12327 8730 12351 8732
rect 12407 8730 12431 8732
rect 12487 8730 12493 8732
rect 12247 8678 12249 8730
rect 12429 8678 12431 8730
rect 12185 8676 12191 8678
rect 12247 8676 12271 8678
rect 12327 8676 12351 8678
rect 12407 8676 12431 8678
rect 12487 8676 12493 8678
rect 12185 8667 12493 8676
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 12544 8430 12572 8978
rect 12636 8906 12664 9658
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12728 8974 12756 9522
rect 12820 9058 12848 10610
rect 13096 10169 13124 11222
rect 13360 11212 13412 11218
rect 13360 11154 13412 11160
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13082 10160 13138 10169
rect 13280 10130 13308 10746
rect 13372 10538 13400 11154
rect 13464 10742 13492 11766
rect 13740 11694 13768 12242
rect 14476 11762 14504 12310
rect 15212 11898 15240 13126
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 14188 11620 14240 11626
rect 14188 11562 14240 11568
rect 14200 11218 14228 11562
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13636 10600 13688 10606
rect 13688 10548 13768 10554
rect 13636 10542 13768 10548
rect 13360 10532 13412 10538
rect 13648 10526 13768 10542
rect 13360 10474 13412 10480
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13082 10095 13138 10104
rect 13176 10124 13228 10130
rect 12900 9988 12952 9994
rect 12900 9930 12952 9936
rect 12912 9178 12940 9930
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9654 13032 9862
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12820 9030 12940 9058
rect 13096 9042 13124 10095
rect 13176 10066 13228 10072
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13188 9586 13216 10066
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13176 9580 13228 9586
rect 13176 9522 13228 9528
rect 13280 9178 13308 9862
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12636 8090 12664 8842
rect 12728 8650 12756 8910
rect 12728 8622 12848 8650
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12728 8090 12756 8366
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12185 7644 12493 7653
rect 12185 7642 12191 7644
rect 12247 7642 12271 7644
rect 12327 7642 12351 7644
rect 12407 7642 12431 7644
rect 12487 7642 12493 7644
rect 12247 7590 12249 7642
rect 12429 7590 12431 7642
rect 12185 7588 12191 7590
rect 12247 7588 12271 7590
rect 12327 7588 12351 7590
rect 12407 7588 12431 7590
rect 12487 7588 12493 7590
rect 12185 7579 12493 7588
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6860 11020 6866
rect 11072 6848 11100 7142
rect 11532 6934 11560 7278
rect 11520 6928 11572 6934
rect 11020 6820 11100 6848
rect 11150 6896 11206 6905
rect 11520 6870 11572 6876
rect 11150 6831 11152 6840
rect 10968 6802 11020 6808
rect 11204 6831 11206 6840
rect 11336 6860 11388 6866
rect 11152 6802 11204 6808
rect 11336 6802 11388 6808
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10324 6248 10376 6254
rect 10324 6190 10376 6196
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10152 5778 10272 5794
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 10140 5772 10272 5778
rect 10192 5766 10272 5772
rect 11060 5772 11112 5778
rect 10140 5714 10192 5720
rect 11060 5714 11112 5720
rect 11072 5234 11100 5714
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 9827 4924 10135 4933
rect 9827 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10073 4924
rect 10129 4922 10135 4924
rect 9889 4870 9891 4922
rect 10071 4870 10073 4922
rect 9827 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10073 4870
rect 10129 4868 10135 4870
rect 9827 4859 10135 4868
rect 9827 3836 10135 3845
rect 9827 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10073 3836
rect 10129 3834 10135 3836
rect 9889 3782 9891 3834
rect 10071 3782 10073 3834
rect 9827 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10073 3782
rect 10129 3780 10135 3782
rect 9827 3771 10135 3780
rect 9827 2748 10135 2757
rect 9827 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10073 2748
rect 10129 2746 10135 2748
rect 9889 2694 9891 2746
rect 10071 2694 10073 2746
rect 9827 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10073 2694
rect 10129 2692 10135 2694
rect 9827 2683 10135 2692
rect 9827 1660 10135 1669
rect 9827 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10073 1660
rect 10129 1658 10135 1660
rect 9889 1606 9891 1658
rect 10071 1606 10073 1658
rect 9827 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10073 1606
rect 10129 1604 10135 1606
rect 9827 1595 10135 1604
rect 9827 572 10135 581
rect 9827 570 9833 572
rect 9889 570 9913 572
rect 9969 570 9993 572
rect 10049 570 10073 572
rect 10129 570 10135 572
rect 9889 518 9891 570
rect 10071 518 10073 570
rect 9827 516 9833 518
rect 9889 516 9913 518
rect 9969 516 9993 518
rect 10049 516 10073 518
rect 10129 516 10135 518
rect 9827 507 10135 516
rect 11164 400 11192 5510
rect 11256 5166 11284 6598
rect 11348 6186 11376 6802
rect 11808 6798 11836 7278
rect 12072 7268 12124 7274
rect 12072 7210 12124 7216
rect 12164 7268 12216 7274
rect 12544 7256 12572 7958
rect 12636 7342 12664 8026
rect 12820 7478 12848 8622
rect 12912 7954 12940 9030
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13188 8634 13216 8978
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13188 8514 13216 8570
rect 13004 8486 13216 8514
rect 13280 8498 13308 9114
rect 13268 8492 13320 8498
rect 12900 7948 12952 7954
rect 12900 7890 12952 7896
rect 12912 7750 12940 7890
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12808 7472 12860 7478
rect 12808 7414 12860 7420
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12216 7228 12572 7256
rect 12164 7210 12216 7216
rect 12084 7002 12112 7210
rect 12636 7002 12664 7278
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 6866 12756 7278
rect 12820 7274 12848 7414
rect 13004 7342 13032 8486
rect 13268 8434 13320 8440
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13188 7954 13216 8366
rect 13556 8090 13584 10406
rect 13634 10296 13690 10305
rect 13634 10231 13636 10240
rect 13688 10231 13690 10240
rect 13636 10202 13688 10208
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13648 10033 13676 10066
rect 13634 10024 13690 10033
rect 13634 9959 13690 9968
rect 13740 9518 13768 10526
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 9042 13768 9454
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13832 8430 13860 11018
rect 14200 10742 14228 11154
rect 14476 11150 14504 11698
rect 15212 11694 15240 11834
rect 15304 11694 15332 14486
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15200 11688 15252 11694
rect 15200 11630 15252 11636
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14542 11452 14850 11461
rect 14542 11450 14548 11452
rect 14604 11450 14628 11452
rect 14684 11450 14708 11452
rect 14764 11450 14788 11452
rect 14844 11450 14850 11452
rect 14604 11398 14606 11450
rect 14786 11398 14788 11450
rect 14542 11396 14548 11398
rect 14604 11396 14628 11398
rect 14684 11396 14708 11398
rect 14764 11396 14788 11398
rect 14844 11396 14850 11398
rect 14542 11387 14850 11396
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 10810 14504 10950
rect 14752 10810 14780 11154
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14740 10804 14792 10810
rect 14740 10746 14792 10752
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14936 10606 14964 11562
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11286 15332 11494
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15108 11212 15160 11218
rect 15028 11172 15108 11200
rect 15028 10742 15056 11172
rect 15108 11154 15160 11160
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 15120 10606 15148 10950
rect 15304 10742 15332 10950
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 13924 10198 13952 10406
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 14016 10062 14044 10406
rect 14200 10266 14228 10542
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 10305 14412 10406
rect 14542 10364 14850 10373
rect 14542 10362 14548 10364
rect 14604 10362 14628 10364
rect 14684 10362 14708 10364
rect 14764 10362 14788 10364
rect 14844 10362 14850 10364
rect 14604 10310 14606 10362
rect 14786 10310 14788 10362
rect 14542 10308 14548 10310
rect 14604 10308 14628 10310
rect 14684 10308 14708 10310
rect 14764 10308 14788 10310
rect 14844 10308 14850 10310
rect 14370 10296 14426 10305
rect 14542 10299 14850 10308
rect 14188 10260 14240 10266
rect 14370 10231 14426 10240
rect 14188 10202 14240 10208
rect 14200 10169 14228 10202
rect 14186 10160 14242 10169
rect 14242 10130 14688 10146
rect 14242 10124 14700 10130
rect 14242 10118 14648 10124
rect 14186 10095 14242 10104
rect 14648 10066 14700 10072
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14738 10024 14794 10033
rect 14384 9722 14412 9998
rect 14738 9959 14740 9968
rect 14792 9959 14794 9968
rect 14740 9930 14792 9936
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14108 9602 14136 9658
rect 13924 9574 14136 9602
rect 14464 9580 14516 9586
rect 13924 9518 13952 9574
rect 14464 9522 14516 9528
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 14108 8294 14136 8570
rect 14476 8430 14504 9522
rect 14542 9276 14850 9285
rect 14542 9274 14548 9276
rect 14604 9274 14628 9276
rect 14684 9274 14708 9276
rect 14764 9274 14788 9276
rect 14844 9274 14850 9276
rect 14604 9222 14606 9274
rect 14786 9222 14788 9274
rect 14542 9220 14548 9222
rect 14604 9220 14628 9222
rect 14684 9220 14708 9222
rect 14764 9220 14788 9222
rect 14844 9220 14850 9222
rect 14542 9211 14850 9220
rect 14936 8498 14964 10542
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15028 8906 15056 10406
rect 15212 10266 15240 10406
rect 15396 10266 15424 11834
rect 15488 11558 15516 14758
rect 16224 13870 16252 14826
rect 19257 14716 19565 14725
rect 19257 14714 19263 14716
rect 19319 14714 19343 14716
rect 19399 14714 19423 14716
rect 19479 14714 19503 14716
rect 19559 14714 19565 14716
rect 19319 14662 19321 14714
rect 19501 14662 19503 14714
rect 19257 14660 19263 14662
rect 19319 14660 19343 14662
rect 19399 14660 19423 14662
rect 19479 14660 19503 14662
rect 19559 14660 19565 14662
rect 19257 14651 19565 14660
rect 16900 14172 17208 14181
rect 16900 14170 16906 14172
rect 16962 14170 16986 14172
rect 17042 14170 17066 14172
rect 17122 14170 17146 14172
rect 17202 14170 17208 14172
rect 16962 14118 16964 14170
rect 17144 14118 17146 14170
rect 16900 14116 16906 14118
rect 16962 14116 16986 14118
rect 17042 14116 17066 14118
rect 17122 14116 17146 14118
rect 17202 14116 17208 14118
rect 16900 14107 17208 14116
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15948 11898 15976 13738
rect 16224 13394 16252 13806
rect 16500 13530 16528 13806
rect 19257 13628 19565 13637
rect 19257 13626 19263 13628
rect 19319 13626 19343 13628
rect 19399 13626 19423 13628
rect 19479 13626 19503 13628
rect 19559 13626 19565 13628
rect 19319 13574 19321 13626
rect 19501 13574 19503 13626
rect 19257 13572 19263 13574
rect 19319 13572 19343 13574
rect 19399 13572 19423 13574
rect 19479 13572 19503 13574
rect 19559 13572 19565 13574
rect 19257 13563 19565 13572
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16500 13394 16528 13466
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 16900 13084 17208 13093
rect 16900 13082 16906 13084
rect 16962 13082 16986 13084
rect 17042 13082 17066 13084
rect 17122 13082 17146 13084
rect 17202 13082 17208 13084
rect 16962 13030 16964 13082
rect 17144 13030 17146 13082
rect 16900 13028 16906 13030
rect 16962 13028 16986 13030
rect 17042 13028 17066 13030
rect 17122 13028 17146 13030
rect 17202 13028 17208 13030
rect 16900 13019 17208 13028
rect 16304 12708 16356 12714
rect 16304 12650 16356 12656
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11218 15516 11494
rect 15764 11218 15792 11698
rect 15948 11506 15976 11834
rect 16316 11694 16344 12650
rect 16900 11996 17208 12005
rect 16900 11994 16906 11996
rect 16962 11994 16986 11996
rect 17042 11994 17066 11996
rect 17122 11994 17146 11996
rect 17202 11994 17208 11996
rect 16962 11942 16964 11994
rect 17144 11942 17146 11994
rect 16900 11940 16906 11942
rect 16962 11940 16986 11942
rect 17042 11940 17066 11942
rect 17122 11940 17146 11942
rect 17202 11940 17208 11942
rect 16900 11931 17208 11940
rect 16672 11824 16724 11830
rect 16672 11766 16724 11772
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 15856 11478 15976 11506
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15212 9518 15240 9658
rect 15396 9586 15424 10202
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15200 9376 15252 9382
rect 15200 9318 15252 9324
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8566 15056 8842
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14936 8378 14964 8434
rect 14096 8288 14148 8294
rect 14096 8230 14148 8236
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13188 7342 13216 7414
rect 13556 7410 13584 7890
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12808 7268 12860 7274
rect 12808 7210 12860 7216
rect 13096 7002 13124 7278
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13464 7002 13492 7210
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13556 6866 13584 7346
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13832 6866 13860 6938
rect 13924 6866 13952 7482
rect 14108 7342 14136 8230
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 6866 14136 7142
rect 14292 7002 14320 7414
rect 14476 7410 14504 8366
rect 14936 8350 15056 8378
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14542 8188 14850 8197
rect 14542 8186 14548 8188
rect 14604 8186 14628 8188
rect 14684 8186 14708 8188
rect 14764 8186 14788 8188
rect 14844 8186 14850 8188
rect 14604 8134 14606 8186
rect 14786 8134 14788 8186
rect 14542 8132 14548 8134
rect 14604 8132 14628 8134
rect 14684 8132 14708 8134
rect 14764 8132 14788 8134
rect 14844 8132 14850 8134
rect 14542 8123 14850 8132
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14844 7546 14872 7822
rect 14936 7818 14964 8230
rect 15028 8022 15056 8350
rect 15016 8016 15068 8022
rect 15016 7958 15068 7964
rect 15212 7818 15240 9318
rect 14924 7812 14976 7818
rect 14924 7754 14976 7760
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 7290 14504 7346
rect 14844 7342 14872 7482
rect 15028 7342 15056 7686
rect 15120 7410 15148 7686
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14384 7262 14504 7290
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 14384 7206 14412 7262
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14280 6996 14332 7002
rect 14280 6938 14332 6944
rect 14292 6866 14320 6938
rect 14476 6866 14504 7142
rect 14542 7100 14850 7109
rect 14542 7098 14548 7100
rect 14604 7098 14628 7100
rect 14684 7098 14708 7100
rect 14764 7098 14788 7100
rect 14844 7098 14850 7100
rect 14604 7046 14606 7098
rect 14786 7046 14788 7098
rect 14542 7044 14548 7046
rect 14604 7044 14628 7046
rect 14684 7044 14708 7046
rect 14764 7044 14788 7046
rect 14844 7044 14850 7046
rect 14542 7035 14850 7044
rect 15304 6866 15332 9318
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15396 8498 15424 8774
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15488 8294 15516 10746
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 7954 15516 8230
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15580 7546 15608 10950
rect 15672 10674 15700 11154
rect 15856 10810 15884 11478
rect 16040 11354 16068 11630
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15856 10606 15884 10746
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 9518 15792 10134
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 9036 15712 9042
rect 15660 8978 15712 8984
rect 15672 8430 15700 8978
rect 15856 8974 15884 10406
rect 15948 9364 15976 11290
rect 16040 11218 16068 11290
rect 16316 11218 16344 11630
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16028 11212 16080 11218
rect 16028 11154 16080 11160
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16316 10674 16344 11154
rect 16408 11082 16436 11494
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16500 11200 16528 11290
rect 16684 11218 16712 11766
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16672 11212 16724 11218
rect 16500 11172 16620 11200
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16408 10674 16436 11018
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16028 10464 16080 10470
rect 16028 10406 16080 10412
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16040 10198 16068 10406
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 15948 9336 16068 9364
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8430 15884 8910
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15752 8424 15804 8430
rect 15752 8366 15804 8372
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15568 7540 15620 7546
rect 15568 7482 15620 7488
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 6934 15608 7142
rect 15672 6934 15700 8366
rect 15764 8090 15792 8366
rect 15948 8090 15976 8978
rect 16040 8430 16068 9336
rect 16132 8838 16160 9998
rect 16224 9450 16252 10066
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9518 16344 9862
rect 16500 9722 16528 10406
rect 16592 9994 16620 11172
rect 16672 11154 16724 11160
rect 16776 10606 16804 11698
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11218 16896 11494
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 17224 11212 17276 11218
rect 17224 11154 17276 11160
rect 16900 10908 17208 10917
rect 16900 10906 16906 10908
rect 16962 10906 16986 10908
rect 17042 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17208 10908
rect 16962 10854 16964 10906
rect 17144 10854 17146 10906
rect 16900 10852 16906 10854
rect 16962 10852 16986 10854
rect 17042 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17208 10854
rect 16900 10843 17208 10852
rect 17236 10742 17264 11154
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16488 9716 16540 9722
rect 16488 9658 16540 9664
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8430 16160 8774
rect 16028 8424 16080 8430
rect 16028 8366 16080 8372
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15764 7834 15792 8026
rect 15764 7806 15884 7834
rect 15856 7342 15884 7806
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15568 6928 15620 6934
rect 15568 6870 15620 6876
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14280 6860 14332 6866
rect 14280 6802 14332 6808
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15292 6860 15344 6866
rect 15292 6802 15344 6808
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 12185 6556 12493 6565
rect 12185 6554 12191 6556
rect 12247 6554 12271 6556
rect 12327 6554 12351 6556
rect 12407 6554 12431 6556
rect 12487 6554 12493 6556
rect 12247 6502 12249 6554
rect 12429 6502 12431 6554
rect 12185 6500 12191 6502
rect 12247 6500 12271 6502
rect 12327 6500 12351 6502
rect 12407 6500 12431 6502
rect 12487 6500 12493 6502
rect 12185 6491 12493 6500
rect 12544 6458 12572 6802
rect 14568 6458 14596 6802
rect 15212 6730 15240 6802
rect 16040 6798 16068 8366
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16316 8090 16344 8230
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16408 7954 16436 8298
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16500 7478 16528 9658
rect 16592 8430 16620 9930
rect 16900 9820 17208 9829
rect 16900 9818 16906 9820
rect 16962 9818 16986 9820
rect 17042 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17208 9820
rect 16962 9766 16964 9818
rect 17144 9766 17146 9818
rect 16900 9764 16906 9766
rect 16962 9764 16986 9766
rect 17042 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17208 9766
rect 16900 9755 17208 9764
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16684 9518 16712 9590
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 8498 16712 9454
rect 17236 9178 17264 10678
rect 17500 10600 17552 10606
rect 17500 10542 17552 10548
rect 17316 10124 17368 10130
rect 17316 10066 17368 10072
rect 17328 9926 17356 10066
rect 17316 9920 17368 9926
rect 17316 9862 17368 9868
rect 17328 9586 17356 9862
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17236 8974 17264 9114
rect 17328 9042 17356 9522
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 16900 8732 17208 8741
rect 16900 8730 16906 8732
rect 16962 8730 16986 8732
rect 17042 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17208 8732
rect 16962 8678 16964 8730
rect 17144 8678 17146 8730
rect 16900 8676 16906 8678
rect 16962 8676 16986 8678
rect 17042 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17208 8678
rect 16900 8667 17208 8676
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16684 7970 16712 8434
rect 16776 8294 16804 8570
rect 17236 8514 17264 8910
rect 17144 8486 17264 8514
rect 17420 8498 17448 8910
rect 17144 8430 17172 8486
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16592 7954 16712 7970
rect 16580 7948 16712 7954
rect 16632 7942 16712 7948
rect 16580 7890 16632 7896
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6798 16436 7142
rect 16500 6866 16528 7414
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11532 5778 11560 6326
rect 14542 6012 14850 6021
rect 14542 6010 14548 6012
rect 14604 6010 14628 6012
rect 14684 6010 14708 6012
rect 14764 6010 14788 6012
rect 14844 6010 14850 6012
rect 14604 5958 14606 6010
rect 14786 5958 14788 6010
rect 14542 5956 14548 5958
rect 14604 5956 14628 5958
rect 14684 5956 14708 5958
rect 14764 5956 14788 5958
rect 14844 5956 14850 5958
rect 14542 5947 14850 5956
rect 16592 5846 16620 7754
rect 16684 7342 16712 7942
rect 16776 7546 16804 8230
rect 16868 7818 16896 8366
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16900 7644 17208 7653
rect 16900 7642 16906 7644
rect 16962 7642 16986 7644
rect 17042 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17208 7644
rect 16962 7590 16964 7642
rect 17144 7590 17146 7642
rect 16900 7588 16906 7590
rect 16962 7588 16986 7590
rect 17042 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17208 7590
rect 16900 7579 17208 7588
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 17236 7410 17264 8486
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17512 8022 17540 10542
rect 17880 10470 17908 13126
rect 19257 12540 19565 12549
rect 19257 12538 19263 12540
rect 19319 12538 19343 12540
rect 19399 12538 19423 12540
rect 19479 12538 19503 12540
rect 19559 12538 19565 12540
rect 19319 12486 19321 12538
rect 19501 12486 19503 12538
rect 19257 12484 19263 12486
rect 19319 12484 19343 12486
rect 19399 12484 19423 12486
rect 19479 12484 19503 12486
rect 19559 12484 19565 12486
rect 19257 12475 19565 12484
rect 19257 11452 19565 11461
rect 19257 11450 19263 11452
rect 19319 11450 19343 11452
rect 19399 11450 19423 11452
rect 19479 11450 19503 11452
rect 19559 11450 19565 11452
rect 19319 11398 19321 11450
rect 19501 11398 19503 11450
rect 19257 11396 19263 11398
rect 19319 11396 19343 11398
rect 19399 11396 19423 11398
rect 19479 11396 19503 11398
rect 19559 11396 19565 11398
rect 19257 11387 19565 11396
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10266 17908 10406
rect 19257 10364 19565 10373
rect 19257 10362 19263 10364
rect 19319 10362 19343 10364
rect 19399 10362 19423 10364
rect 19479 10362 19503 10364
rect 19559 10362 19565 10364
rect 19319 10310 19321 10362
rect 19501 10310 19503 10362
rect 19257 10308 19263 10310
rect 19319 10308 19343 10310
rect 19399 10308 19423 10310
rect 19479 10308 19503 10310
rect 19559 10308 19565 10310
rect 19257 10299 19565 10308
rect 17868 10260 17920 10266
rect 17868 10202 17920 10208
rect 17880 10010 17908 10202
rect 17880 9982 18092 10010
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 8514 17908 9862
rect 17880 8498 18000 8514
rect 17880 8492 18012 8498
rect 17880 8486 17960 8492
rect 17960 8434 18012 8440
rect 18064 8362 18092 9982
rect 19257 9276 19565 9285
rect 19257 9274 19263 9276
rect 19319 9274 19343 9276
rect 19399 9274 19423 9276
rect 19479 9274 19503 9276
rect 19559 9274 19565 9276
rect 19319 9222 19321 9274
rect 19501 9222 19503 9274
rect 19257 9220 19263 9222
rect 19319 9220 19343 9222
rect 19399 9220 19423 9222
rect 19479 9220 19503 9222
rect 19559 9220 19565 9222
rect 19257 9211 19565 9220
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 8634 18368 8978
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17880 7954 17908 8230
rect 19257 8188 19565 8197
rect 19257 8186 19263 8188
rect 19319 8186 19343 8188
rect 19399 8186 19423 8188
rect 19479 8186 19503 8188
rect 19559 8186 19565 8188
rect 19319 8134 19321 8186
rect 19501 8134 19503 8186
rect 19257 8132 19263 8134
rect 19319 8132 19343 8134
rect 19399 8132 19423 8134
rect 19479 8132 19503 8134
rect 19559 8132 19565 8134
rect 19257 8123 19565 8132
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 19257 7100 19565 7109
rect 19257 7098 19263 7100
rect 19319 7098 19343 7100
rect 19399 7098 19423 7100
rect 19479 7098 19503 7100
rect 19559 7098 19565 7100
rect 19319 7046 19321 7098
rect 19501 7046 19503 7098
rect 19257 7044 19263 7046
rect 19319 7044 19343 7046
rect 19399 7044 19423 7046
rect 19479 7044 19503 7046
rect 19559 7044 19565 7046
rect 19257 7035 19565 7044
rect 16900 6556 17208 6565
rect 16900 6554 16906 6556
rect 16962 6554 16986 6556
rect 17042 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17208 6556
rect 16962 6502 16964 6554
rect 17144 6502 17146 6554
rect 16900 6500 16906 6502
rect 16962 6500 16986 6502
rect 17042 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17208 6502
rect 16900 6491 17208 6500
rect 19257 6012 19565 6021
rect 19257 6010 19263 6012
rect 19319 6010 19343 6012
rect 19399 6010 19423 6012
rect 19479 6010 19503 6012
rect 19559 6010 19565 6012
rect 19319 5958 19321 6010
rect 19501 5958 19503 6010
rect 19257 5956 19263 5958
rect 19319 5956 19343 5958
rect 19399 5956 19423 5958
rect 19479 5956 19503 5958
rect 19559 5956 19565 5958
rect 19257 5947 19565 5956
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 18604 5568 18656 5574
rect 18604 5510 18656 5516
rect 12185 5468 12493 5477
rect 12185 5466 12191 5468
rect 12247 5466 12271 5468
rect 12327 5466 12351 5468
rect 12407 5466 12431 5468
rect 12487 5466 12493 5468
rect 12247 5414 12249 5466
rect 12429 5414 12431 5466
rect 12185 5412 12191 5414
rect 12247 5412 12271 5414
rect 12327 5412 12351 5414
rect 12407 5412 12431 5414
rect 12487 5412 12493 5414
rect 12185 5403 12493 5412
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 12185 4380 12493 4389
rect 12185 4378 12191 4380
rect 12247 4378 12271 4380
rect 12327 4378 12351 4380
rect 12407 4378 12431 4380
rect 12487 4378 12493 4380
rect 12247 4326 12249 4378
rect 12429 4326 12431 4378
rect 12185 4324 12191 4326
rect 12247 4324 12271 4326
rect 12327 4324 12351 4326
rect 12407 4324 12431 4326
rect 12487 4324 12493 4326
rect 12185 4315 12493 4324
rect 12185 3292 12493 3301
rect 12185 3290 12191 3292
rect 12247 3290 12271 3292
rect 12327 3290 12351 3292
rect 12407 3290 12431 3292
rect 12487 3290 12493 3292
rect 12247 3238 12249 3290
rect 12429 3238 12431 3290
rect 12185 3236 12191 3238
rect 12247 3236 12271 3238
rect 12327 3236 12351 3238
rect 12407 3236 12431 3238
rect 12487 3236 12493 3238
rect 12185 3227 12493 3236
rect 12185 2204 12493 2213
rect 12185 2202 12191 2204
rect 12247 2202 12271 2204
rect 12327 2202 12351 2204
rect 12407 2202 12431 2204
rect 12487 2202 12493 2204
rect 12247 2150 12249 2202
rect 12429 2150 12431 2202
rect 12185 2148 12191 2150
rect 12247 2148 12271 2150
rect 12327 2148 12351 2150
rect 12407 2148 12431 2150
rect 12487 2148 12493 2150
rect 12185 2139 12493 2148
rect 12185 1116 12493 1125
rect 12185 1114 12191 1116
rect 12247 1114 12271 1116
rect 12327 1114 12351 1116
rect 12407 1114 12431 1116
rect 12487 1114 12493 1116
rect 12247 1062 12249 1114
rect 12429 1062 12431 1114
rect 12185 1060 12191 1062
rect 12247 1060 12271 1062
rect 12327 1060 12351 1062
rect 12407 1060 12431 1062
rect 12487 1060 12493 1062
rect 12185 1051 12493 1060
rect 13648 400 13676 4966
rect 14542 4924 14850 4933
rect 14542 4922 14548 4924
rect 14604 4922 14628 4924
rect 14684 4922 14708 4924
rect 14764 4922 14788 4924
rect 14844 4922 14850 4924
rect 14604 4870 14606 4922
rect 14786 4870 14788 4922
rect 14542 4868 14548 4870
rect 14604 4868 14628 4870
rect 14684 4868 14708 4870
rect 14764 4868 14788 4870
rect 14844 4868 14850 4870
rect 14542 4859 14850 4868
rect 14542 3836 14850 3845
rect 14542 3834 14548 3836
rect 14604 3834 14628 3836
rect 14684 3834 14708 3836
rect 14764 3834 14788 3836
rect 14844 3834 14850 3836
rect 14604 3782 14606 3834
rect 14786 3782 14788 3834
rect 14542 3780 14548 3782
rect 14604 3780 14628 3782
rect 14684 3780 14708 3782
rect 14764 3780 14788 3782
rect 14844 3780 14850 3782
rect 14542 3771 14850 3780
rect 14542 2748 14850 2757
rect 14542 2746 14548 2748
rect 14604 2746 14628 2748
rect 14684 2746 14708 2748
rect 14764 2746 14788 2748
rect 14844 2746 14850 2748
rect 14604 2694 14606 2746
rect 14786 2694 14788 2746
rect 14542 2692 14548 2694
rect 14604 2692 14628 2694
rect 14684 2692 14708 2694
rect 14764 2692 14788 2694
rect 14844 2692 14850 2694
rect 14542 2683 14850 2692
rect 14542 1660 14850 1669
rect 14542 1658 14548 1660
rect 14604 1658 14628 1660
rect 14684 1658 14708 1660
rect 14764 1658 14788 1660
rect 14844 1658 14850 1660
rect 14604 1606 14606 1658
rect 14786 1606 14788 1658
rect 14542 1604 14548 1606
rect 14604 1604 14628 1606
rect 14684 1604 14708 1606
rect 14764 1604 14788 1606
rect 14844 1604 14850 1606
rect 14542 1595 14850 1604
rect 14542 572 14850 581
rect 14542 570 14548 572
rect 14604 570 14628 572
rect 14684 570 14708 572
rect 14764 570 14788 572
rect 14844 570 14850 572
rect 14604 518 14606 570
rect 14786 518 14788 570
rect 14542 516 14548 518
rect 14604 516 14628 518
rect 14684 516 14708 518
rect 14764 516 14788 518
rect 14844 516 14850 518
rect 14542 507 14850 516
rect 16132 400 16160 5510
rect 16900 5468 17208 5477
rect 16900 5466 16906 5468
rect 16962 5466 16986 5468
rect 17042 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17208 5468
rect 16962 5414 16964 5466
rect 17144 5414 17146 5466
rect 16900 5412 16906 5414
rect 16962 5412 16986 5414
rect 17042 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17208 5414
rect 16900 5403 17208 5412
rect 16900 4380 17208 4389
rect 16900 4378 16906 4380
rect 16962 4378 16986 4380
rect 17042 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17208 4380
rect 16962 4326 16964 4378
rect 17144 4326 17146 4378
rect 16900 4324 16906 4326
rect 16962 4324 16986 4326
rect 17042 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17208 4326
rect 16900 4315 17208 4324
rect 16900 3292 17208 3301
rect 16900 3290 16906 3292
rect 16962 3290 16986 3292
rect 17042 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17208 3292
rect 16962 3238 16964 3290
rect 17144 3238 17146 3290
rect 16900 3236 16906 3238
rect 16962 3236 16986 3238
rect 17042 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17208 3238
rect 16900 3227 17208 3236
rect 16900 2204 17208 2213
rect 16900 2202 16906 2204
rect 16962 2202 16986 2204
rect 17042 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17208 2204
rect 16962 2150 16964 2202
rect 17144 2150 17146 2202
rect 16900 2148 16906 2150
rect 16962 2148 16986 2150
rect 17042 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17208 2150
rect 16900 2139 17208 2148
rect 16900 1116 17208 1125
rect 16900 1114 16906 1116
rect 16962 1114 16986 1116
rect 17042 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17208 1116
rect 16962 1062 16964 1114
rect 17144 1062 17146 1114
rect 16900 1060 16906 1062
rect 16962 1060 16986 1062
rect 17042 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17208 1062
rect 16900 1051 17208 1060
rect 18616 400 18644 5510
rect 19257 4924 19565 4933
rect 19257 4922 19263 4924
rect 19319 4922 19343 4924
rect 19399 4922 19423 4924
rect 19479 4922 19503 4924
rect 19559 4922 19565 4924
rect 19319 4870 19321 4922
rect 19501 4870 19503 4922
rect 19257 4868 19263 4870
rect 19319 4868 19343 4870
rect 19399 4868 19423 4870
rect 19479 4868 19503 4870
rect 19559 4868 19565 4870
rect 19257 4859 19565 4868
rect 19257 3836 19565 3845
rect 19257 3834 19263 3836
rect 19319 3834 19343 3836
rect 19399 3834 19423 3836
rect 19479 3834 19503 3836
rect 19559 3834 19565 3836
rect 19319 3782 19321 3834
rect 19501 3782 19503 3834
rect 19257 3780 19263 3782
rect 19319 3780 19343 3782
rect 19399 3780 19423 3782
rect 19479 3780 19503 3782
rect 19559 3780 19565 3782
rect 19257 3771 19565 3780
rect 19257 2748 19565 2757
rect 19257 2746 19263 2748
rect 19319 2746 19343 2748
rect 19399 2746 19423 2748
rect 19479 2746 19503 2748
rect 19559 2746 19565 2748
rect 19319 2694 19321 2746
rect 19501 2694 19503 2746
rect 19257 2692 19263 2694
rect 19319 2692 19343 2694
rect 19399 2692 19423 2694
rect 19479 2692 19503 2694
rect 19559 2692 19565 2694
rect 19257 2683 19565 2692
rect 19257 1660 19565 1669
rect 19257 1658 19263 1660
rect 19319 1658 19343 1660
rect 19399 1658 19423 1660
rect 19479 1658 19503 1660
rect 19559 1658 19565 1660
rect 19319 1606 19321 1658
rect 19501 1606 19503 1658
rect 19257 1604 19263 1606
rect 19319 1604 19343 1606
rect 19399 1604 19423 1606
rect 19479 1604 19503 1606
rect 19559 1604 19565 1606
rect 19257 1595 19565 1604
rect 19257 572 19565 581
rect 19257 570 19263 572
rect 19319 570 19343 572
rect 19399 570 19423 572
rect 19479 570 19503 572
rect 19559 570 19565 572
rect 19319 518 19321 570
rect 19501 518 19503 570
rect 19257 516 19263 518
rect 19319 516 19343 518
rect 19399 516 19423 518
rect 19479 516 19503 518
rect 19559 516 19565 518
rect 19257 507 19565 516
rect 1214 0 1270 400
rect 3698 0 3754 400
rect 6182 0 6238 400
rect 8666 0 8722 400
rect 11150 0 11206 400
rect 13634 0 13690 400
rect 16118 0 16174 400
rect 18602 0 18658 400
<< via2 >>
rect 5118 19066 5174 19068
rect 5198 19066 5254 19068
rect 5278 19066 5334 19068
rect 5358 19066 5414 19068
rect 5118 19014 5164 19066
rect 5164 19014 5174 19066
rect 5198 19014 5228 19066
rect 5228 19014 5240 19066
rect 5240 19014 5254 19066
rect 5278 19014 5292 19066
rect 5292 19014 5304 19066
rect 5304 19014 5334 19066
rect 5358 19014 5368 19066
rect 5368 19014 5414 19066
rect 5118 19012 5174 19014
rect 5198 19012 5254 19014
rect 5278 19012 5334 19014
rect 5358 19012 5414 19014
rect 2761 18522 2817 18524
rect 2841 18522 2897 18524
rect 2921 18522 2977 18524
rect 3001 18522 3057 18524
rect 2761 18470 2807 18522
rect 2807 18470 2817 18522
rect 2841 18470 2871 18522
rect 2871 18470 2883 18522
rect 2883 18470 2897 18522
rect 2921 18470 2935 18522
rect 2935 18470 2947 18522
rect 2947 18470 2977 18522
rect 3001 18470 3011 18522
rect 3011 18470 3057 18522
rect 2761 18468 2817 18470
rect 2841 18468 2897 18470
rect 2921 18468 2977 18470
rect 3001 18468 3057 18470
rect 2761 17434 2817 17436
rect 2841 17434 2897 17436
rect 2921 17434 2977 17436
rect 3001 17434 3057 17436
rect 2761 17382 2807 17434
rect 2807 17382 2817 17434
rect 2841 17382 2871 17434
rect 2871 17382 2883 17434
rect 2883 17382 2897 17434
rect 2921 17382 2935 17434
rect 2935 17382 2947 17434
rect 2947 17382 2977 17434
rect 3001 17382 3011 17434
rect 3011 17382 3057 17434
rect 2761 17380 2817 17382
rect 2841 17380 2897 17382
rect 2921 17380 2977 17382
rect 3001 17380 3057 17382
rect 2761 16346 2817 16348
rect 2841 16346 2897 16348
rect 2921 16346 2977 16348
rect 3001 16346 3057 16348
rect 2761 16294 2807 16346
rect 2807 16294 2817 16346
rect 2841 16294 2871 16346
rect 2871 16294 2883 16346
rect 2883 16294 2897 16346
rect 2921 16294 2935 16346
rect 2935 16294 2947 16346
rect 2947 16294 2977 16346
rect 3001 16294 3011 16346
rect 3011 16294 3057 16346
rect 2761 16292 2817 16294
rect 2841 16292 2897 16294
rect 2921 16292 2977 16294
rect 3001 16292 3057 16294
rect 2761 15258 2817 15260
rect 2841 15258 2897 15260
rect 2921 15258 2977 15260
rect 3001 15258 3057 15260
rect 2761 15206 2807 15258
rect 2807 15206 2817 15258
rect 2841 15206 2871 15258
rect 2871 15206 2883 15258
rect 2883 15206 2897 15258
rect 2921 15206 2935 15258
rect 2935 15206 2947 15258
rect 2947 15206 2977 15258
rect 3001 15206 3011 15258
rect 3011 15206 3057 15258
rect 2761 15204 2817 15206
rect 2841 15204 2897 15206
rect 2921 15204 2977 15206
rect 3001 15204 3057 15206
rect 2761 14170 2817 14172
rect 2841 14170 2897 14172
rect 2921 14170 2977 14172
rect 3001 14170 3057 14172
rect 2761 14118 2807 14170
rect 2807 14118 2817 14170
rect 2841 14118 2871 14170
rect 2871 14118 2883 14170
rect 2883 14118 2897 14170
rect 2921 14118 2935 14170
rect 2935 14118 2947 14170
rect 2947 14118 2977 14170
rect 3001 14118 3011 14170
rect 3011 14118 3057 14170
rect 2761 14116 2817 14118
rect 2841 14116 2897 14118
rect 2921 14116 2977 14118
rect 3001 14116 3057 14118
rect 2761 13082 2817 13084
rect 2841 13082 2897 13084
rect 2921 13082 2977 13084
rect 3001 13082 3057 13084
rect 2761 13030 2807 13082
rect 2807 13030 2817 13082
rect 2841 13030 2871 13082
rect 2871 13030 2883 13082
rect 2883 13030 2897 13082
rect 2921 13030 2935 13082
rect 2935 13030 2947 13082
rect 2947 13030 2977 13082
rect 3001 13030 3011 13082
rect 3011 13030 3057 13082
rect 2761 13028 2817 13030
rect 2841 13028 2897 13030
rect 2921 13028 2977 13030
rect 3001 13028 3057 13030
rect 5118 17978 5174 17980
rect 5198 17978 5254 17980
rect 5278 17978 5334 17980
rect 5358 17978 5414 17980
rect 5118 17926 5164 17978
rect 5164 17926 5174 17978
rect 5198 17926 5228 17978
rect 5228 17926 5240 17978
rect 5240 17926 5254 17978
rect 5278 17926 5292 17978
rect 5292 17926 5304 17978
rect 5304 17926 5334 17978
rect 5358 17926 5368 17978
rect 5368 17926 5414 17978
rect 5118 17924 5174 17926
rect 5198 17924 5254 17926
rect 5278 17924 5334 17926
rect 5358 17924 5414 17926
rect 7476 18522 7532 18524
rect 7556 18522 7612 18524
rect 7636 18522 7692 18524
rect 7716 18522 7772 18524
rect 7476 18470 7522 18522
rect 7522 18470 7532 18522
rect 7556 18470 7586 18522
rect 7586 18470 7598 18522
rect 7598 18470 7612 18522
rect 7636 18470 7650 18522
rect 7650 18470 7662 18522
rect 7662 18470 7692 18522
rect 7716 18470 7726 18522
rect 7726 18470 7772 18522
rect 7476 18468 7532 18470
rect 7556 18468 7612 18470
rect 7636 18468 7692 18470
rect 7716 18468 7772 18470
rect 5118 16890 5174 16892
rect 5198 16890 5254 16892
rect 5278 16890 5334 16892
rect 5358 16890 5414 16892
rect 5118 16838 5164 16890
rect 5164 16838 5174 16890
rect 5198 16838 5228 16890
rect 5228 16838 5240 16890
rect 5240 16838 5254 16890
rect 5278 16838 5292 16890
rect 5292 16838 5304 16890
rect 5304 16838 5334 16890
rect 5358 16838 5368 16890
rect 5368 16838 5414 16890
rect 5118 16836 5174 16838
rect 5198 16836 5254 16838
rect 5278 16836 5334 16838
rect 5358 16836 5414 16838
rect 6182 16668 6184 16688
rect 6184 16668 6236 16688
rect 6236 16668 6238 16688
rect 5118 15802 5174 15804
rect 5198 15802 5254 15804
rect 5278 15802 5334 15804
rect 5358 15802 5414 15804
rect 5118 15750 5164 15802
rect 5164 15750 5174 15802
rect 5198 15750 5228 15802
rect 5228 15750 5240 15802
rect 5240 15750 5254 15802
rect 5278 15750 5292 15802
rect 5292 15750 5304 15802
rect 5304 15750 5334 15802
rect 5358 15750 5368 15802
rect 5368 15750 5414 15802
rect 5118 15748 5174 15750
rect 5198 15748 5254 15750
rect 5278 15748 5334 15750
rect 5358 15748 5414 15750
rect 6182 16632 6238 16668
rect 5118 14714 5174 14716
rect 5198 14714 5254 14716
rect 5278 14714 5334 14716
rect 5358 14714 5414 14716
rect 5118 14662 5164 14714
rect 5164 14662 5174 14714
rect 5198 14662 5228 14714
rect 5228 14662 5240 14714
rect 5240 14662 5254 14714
rect 5278 14662 5292 14714
rect 5292 14662 5304 14714
rect 5304 14662 5334 14714
rect 5358 14662 5368 14714
rect 5368 14662 5414 14714
rect 5118 14660 5174 14662
rect 5198 14660 5254 14662
rect 5278 14660 5334 14662
rect 5358 14660 5414 14662
rect 5118 13626 5174 13628
rect 5198 13626 5254 13628
rect 5278 13626 5334 13628
rect 5358 13626 5414 13628
rect 5118 13574 5164 13626
rect 5164 13574 5174 13626
rect 5198 13574 5228 13626
rect 5228 13574 5240 13626
rect 5240 13574 5254 13626
rect 5278 13574 5292 13626
rect 5292 13574 5304 13626
rect 5304 13574 5334 13626
rect 5358 13574 5368 13626
rect 5368 13574 5414 13626
rect 5118 13572 5174 13574
rect 5198 13572 5254 13574
rect 5278 13572 5334 13574
rect 5358 13572 5414 13574
rect 2761 11994 2817 11996
rect 2841 11994 2897 11996
rect 2921 11994 2977 11996
rect 3001 11994 3057 11996
rect 2761 11942 2807 11994
rect 2807 11942 2817 11994
rect 2841 11942 2871 11994
rect 2871 11942 2883 11994
rect 2883 11942 2897 11994
rect 2921 11942 2935 11994
rect 2935 11942 2947 11994
rect 2947 11942 2977 11994
rect 3001 11942 3011 11994
rect 3011 11942 3057 11994
rect 2761 11940 2817 11942
rect 2841 11940 2897 11942
rect 2921 11940 2977 11942
rect 3001 11940 3057 11942
rect 2761 10906 2817 10908
rect 2841 10906 2897 10908
rect 2921 10906 2977 10908
rect 3001 10906 3057 10908
rect 2761 10854 2807 10906
rect 2807 10854 2817 10906
rect 2841 10854 2871 10906
rect 2871 10854 2883 10906
rect 2883 10854 2897 10906
rect 2921 10854 2935 10906
rect 2935 10854 2947 10906
rect 2947 10854 2977 10906
rect 3001 10854 3011 10906
rect 3011 10854 3057 10906
rect 2761 10852 2817 10854
rect 2841 10852 2897 10854
rect 2921 10852 2977 10854
rect 3001 10852 3057 10854
rect 5118 12538 5174 12540
rect 5198 12538 5254 12540
rect 5278 12538 5334 12540
rect 5358 12538 5414 12540
rect 5118 12486 5164 12538
rect 5164 12486 5174 12538
rect 5198 12486 5228 12538
rect 5228 12486 5240 12538
rect 5240 12486 5254 12538
rect 5278 12486 5292 12538
rect 5292 12486 5304 12538
rect 5304 12486 5334 12538
rect 5358 12486 5368 12538
rect 5368 12486 5414 12538
rect 5118 12484 5174 12486
rect 5198 12484 5254 12486
rect 5278 12484 5334 12486
rect 5358 12484 5414 12486
rect 6918 12724 6920 12744
rect 6920 12724 6972 12744
rect 6972 12724 6974 12744
rect 6918 12688 6974 12724
rect 5118 11450 5174 11452
rect 5198 11450 5254 11452
rect 5278 11450 5334 11452
rect 5358 11450 5414 11452
rect 5118 11398 5164 11450
rect 5164 11398 5174 11450
rect 5198 11398 5228 11450
rect 5228 11398 5240 11450
rect 5240 11398 5254 11450
rect 5278 11398 5292 11450
rect 5292 11398 5304 11450
rect 5304 11398 5334 11450
rect 5358 11398 5368 11450
rect 5368 11398 5414 11450
rect 5118 11396 5174 11398
rect 5198 11396 5254 11398
rect 5278 11396 5334 11398
rect 5358 11396 5414 11398
rect 5118 10362 5174 10364
rect 5198 10362 5254 10364
rect 5278 10362 5334 10364
rect 5358 10362 5414 10364
rect 5118 10310 5164 10362
rect 5164 10310 5174 10362
rect 5198 10310 5228 10362
rect 5228 10310 5240 10362
rect 5240 10310 5254 10362
rect 5278 10310 5292 10362
rect 5292 10310 5304 10362
rect 5304 10310 5334 10362
rect 5358 10310 5368 10362
rect 5368 10310 5414 10362
rect 5118 10308 5174 10310
rect 5198 10308 5254 10310
rect 5278 10308 5334 10310
rect 5358 10308 5414 10310
rect 7476 17434 7532 17436
rect 7556 17434 7612 17436
rect 7636 17434 7692 17436
rect 7716 17434 7772 17436
rect 7476 17382 7522 17434
rect 7522 17382 7532 17434
rect 7556 17382 7586 17434
rect 7586 17382 7598 17434
rect 7598 17382 7612 17434
rect 7636 17382 7650 17434
rect 7650 17382 7662 17434
rect 7662 17382 7692 17434
rect 7716 17382 7726 17434
rect 7726 17382 7772 17434
rect 7476 17380 7532 17382
rect 7556 17380 7612 17382
rect 7636 17380 7692 17382
rect 7716 17380 7772 17382
rect 7476 16346 7532 16348
rect 7556 16346 7612 16348
rect 7636 16346 7692 16348
rect 7716 16346 7772 16348
rect 7476 16294 7522 16346
rect 7522 16294 7532 16346
rect 7556 16294 7586 16346
rect 7586 16294 7598 16346
rect 7598 16294 7612 16346
rect 7636 16294 7650 16346
rect 7650 16294 7662 16346
rect 7662 16294 7692 16346
rect 7716 16294 7726 16346
rect 7726 16294 7772 16346
rect 7476 16292 7532 16294
rect 7556 16292 7612 16294
rect 7636 16292 7692 16294
rect 7716 16292 7772 16294
rect 7476 15258 7532 15260
rect 7556 15258 7612 15260
rect 7636 15258 7692 15260
rect 7716 15258 7772 15260
rect 7476 15206 7522 15258
rect 7522 15206 7532 15258
rect 7556 15206 7586 15258
rect 7586 15206 7598 15258
rect 7598 15206 7612 15258
rect 7636 15206 7650 15258
rect 7650 15206 7662 15258
rect 7662 15206 7692 15258
rect 7716 15206 7726 15258
rect 7726 15206 7772 15258
rect 7476 15204 7532 15206
rect 7556 15204 7612 15206
rect 7636 15204 7692 15206
rect 7716 15204 7772 15206
rect 7476 14170 7532 14172
rect 7556 14170 7612 14172
rect 7636 14170 7692 14172
rect 7716 14170 7772 14172
rect 7476 14118 7522 14170
rect 7522 14118 7532 14170
rect 7556 14118 7586 14170
rect 7586 14118 7598 14170
rect 7598 14118 7612 14170
rect 7636 14118 7650 14170
rect 7650 14118 7662 14170
rect 7662 14118 7692 14170
rect 7716 14118 7726 14170
rect 7726 14118 7772 14170
rect 7476 14116 7532 14118
rect 7556 14116 7612 14118
rect 7636 14116 7692 14118
rect 7716 14116 7772 14118
rect 7476 13082 7532 13084
rect 7556 13082 7612 13084
rect 7636 13082 7692 13084
rect 7716 13082 7772 13084
rect 7476 13030 7522 13082
rect 7522 13030 7532 13082
rect 7556 13030 7586 13082
rect 7586 13030 7598 13082
rect 7598 13030 7612 13082
rect 7636 13030 7650 13082
rect 7650 13030 7662 13082
rect 7662 13030 7692 13082
rect 7716 13030 7726 13082
rect 7726 13030 7772 13082
rect 7476 13028 7532 13030
rect 7556 13028 7612 13030
rect 7636 13028 7692 13030
rect 7716 13028 7772 13030
rect 7476 11994 7532 11996
rect 7556 11994 7612 11996
rect 7636 11994 7692 11996
rect 7716 11994 7772 11996
rect 7476 11942 7522 11994
rect 7522 11942 7532 11994
rect 7556 11942 7586 11994
rect 7586 11942 7598 11994
rect 7598 11942 7612 11994
rect 7636 11942 7650 11994
rect 7650 11942 7662 11994
rect 7662 11942 7692 11994
rect 7716 11942 7726 11994
rect 7726 11942 7772 11994
rect 7476 11940 7532 11942
rect 7556 11940 7612 11942
rect 7636 11940 7692 11942
rect 7716 11940 7772 11942
rect 7476 10906 7532 10908
rect 7556 10906 7612 10908
rect 7636 10906 7692 10908
rect 7716 10906 7772 10908
rect 7476 10854 7522 10906
rect 7522 10854 7532 10906
rect 7556 10854 7586 10906
rect 7586 10854 7598 10906
rect 7598 10854 7612 10906
rect 7636 10854 7650 10906
rect 7650 10854 7662 10906
rect 7662 10854 7692 10906
rect 7716 10854 7726 10906
rect 7726 10854 7772 10906
rect 7476 10852 7532 10854
rect 7556 10852 7612 10854
rect 7636 10852 7692 10854
rect 7716 10852 7772 10854
rect 2761 9818 2817 9820
rect 2841 9818 2897 9820
rect 2921 9818 2977 9820
rect 3001 9818 3057 9820
rect 2761 9766 2807 9818
rect 2807 9766 2817 9818
rect 2841 9766 2871 9818
rect 2871 9766 2883 9818
rect 2883 9766 2897 9818
rect 2921 9766 2935 9818
rect 2935 9766 2947 9818
rect 2947 9766 2977 9818
rect 3001 9766 3011 9818
rect 3011 9766 3057 9818
rect 2761 9764 2817 9766
rect 2841 9764 2897 9766
rect 2921 9764 2977 9766
rect 3001 9764 3057 9766
rect 5118 9274 5174 9276
rect 5198 9274 5254 9276
rect 5278 9274 5334 9276
rect 5358 9274 5414 9276
rect 5118 9222 5164 9274
rect 5164 9222 5174 9274
rect 5198 9222 5228 9274
rect 5228 9222 5240 9274
rect 5240 9222 5254 9274
rect 5278 9222 5292 9274
rect 5292 9222 5304 9274
rect 5304 9222 5334 9274
rect 5358 9222 5368 9274
rect 5368 9222 5414 9274
rect 5118 9220 5174 9222
rect 5198 9220 5254 9222
rect 5278 9220 5334 9222
rect 5358 9220 5414 9222
rect 2761 8730 2817 8732
rect 2841 8730 2897 8732
rect 2921 8730 2977 8732
rect 3001 8730 3057 8732
rect 2761 8678 2807 8730
rect 2807 8678 2817 8730
rect 2841 8678 2871 8730
rect 2871 8678 2883 8730
rect 2883 8678 2897 8730
rect 2921 8678 2935 8730
rect 2935 8678 2947 8730
rect 2947 8678 2977 8730
rect 3001 8678 3011 8730
rect 3011 8678 3057 8730
rect 2761 8676 2817 8678
rect 2841 8676 2897 8678
rect 2921 8676 2977 8678
rect 3001 8676 3057 8678
rect 5118 8186 5174 8188
rect 5198 8186 5254 8188
rect 5278 8186 5334 8188
rect 5358 8186 5414 8188
rect 5118 8134 5164 8186
rect 5164 8134 5174 8186
rect 5198 8134 5228 8186
rect 5228 8134 5240 8186
rect 5240 8134 5254 8186
rect 5278 8134 5292 8186
rect 5292 8134 5304 8186
rect 5304 8134 5334 8186
rect 5358 8134 5368 8186
rect 5368 8134 5414 8186
rect 5118 8132 5174 8134
rect 5198 8132 5254 8134
rect 5278 8132 5334 8134
rect 5358 8132 5414 8134
rect 2761 7642 2817 7644
rect 2841 7642 2897 7644
rect 2921 7642 2977 7644
rect 3001 7642 3057 7644
rect 2761 7590 2807 7642
rect 2807 7590 2817 7642
rect 2841 7590 2871 7642
rect 2871 7590 2883 7642
rect 2883 7590 2897 7642
rect 2921 7590 2935 7642
rect 2935 7590 2947 7642
rect 2947 7590 2977 7642
rect 3001 7590 3011 7642
rect 3011 7590 3057 7642
rect 2761 7588 2817 7590
rect 2841 7588 2897 7590
rect 2921 7588 2977 7590
rect 3001 7588 3057 7590
rect 5118 7098 5174 7100
rect 5198 7098 5254 7100
rect 5278 7098 5334 7100
rect 5358 7098 5414 7100
rect 5118 7046 5164 7098
rect 5164 7046 5174 7098
rect 5198 7046 5228 7098
rect 5228 7046 5240 7098
rect 5240 7046 5254 7098
rect 5278 7046 5292 7098
rect 5292 7046 5304 7098
rect 5304 7046 5334 7098
rect 5358 7046 5368 7098
rect 5368 7046 5414 7098
rect 5118 7044 5174 7046
rect 5198 7044 5254 7046
rect 5278 7044 5334 7046
rect 5358 7044 5414 7046
rect 2761 6554 2817 6556
rect 2841 6554 2897 6556
rect 2921 6554 2977 6556
rect 3001 6554 3057 6556
rect 2761 6502 2807 6554
rect 2807 6502 2817 6554
rect 2841 6502 2871 6554
rect 2871 6502 2883 6554
rect 2883 6502 2897 6554
rect 2921 6502 2935 6554
rect 2935 6502 2947 6554
rect 2947 6502 2977 6554
rect 3001 6502 3011 6554
rect 3011 6502 3057 6554
rect 2761 6500 2817 6502
rect 2841 6500 2897 6502
rect 2921 6500 2977 6502
rect 3001 6500 3057 6502
rect 5118 6010 5174 6012
rect 5198 6010 5254 6012
rect 5278 6010 5334 6012
rect 5358 6010 5414 6012
rect 5118 5958 5164 6010
rect 5164 5958 5174 6010
rect 5198 5958 5228 6010
rect 5228 5958 5240 6010
rect 5240 5958 5254 6010
rect 5278 5958 5292 6010
rect 5292 5958 5304 6010
rect 5304 5958 5334 6010
rect 5358 5958 5368 6010
rect 5368 5958 5414 6010
rect 5118 5956 5174 5958
rect 5198 5956 5254 5958
rect 5278 5956 5334 5958
rect 5358 5956 5414 5958
rect 2761 5466 2817 5468
rect 2841 5466 2897 5468
rect 2921 5466 2977 5468
rect 3001 5466 3057 5468
rect 2761 5414 2807 5466
rect 2807 5414 2817 5466
rect 2841 5414 2871 5466
rect 2871 5414 2883 5466
rect 2883 5414 2897 5466
rect 2921 5414 2935 5466
rect 2935 5414 2947 5466
rect 2947 5414 2977 5466
rect 3001 5414 3011 5466
rect 3011 5414 3057 5466
rect 2761 5412 2817 5414
rect 2841 5412 2897 5414
rect 2921 5412 2977 5414
rect 3001 5412 3057 5414
rect 5118 4922 5174 4924
rect 5198 4922 5254 4924
rect 5278 4922 5334 4924
rect 5358 4922 5414 4924
rect 5118 4870 5164 4922
rect 5164 4870 5174 4922
rect 5198 4870 5228 4922
rect 5228 4870 5240 4922
rect 5240 4870 5254 4922
rect 5278 4870 5292 4922
rect 5292 4870 5304 4922
rect 5304 4870 5334 4922
rect 5358 4870 5368 4922
rect 5368 4870 5414 4922
rect 5118 4868 5174 4870
rect 5198 4868 5254 4870
rect 5278 4868 5334 4870
rect 5358 4868 5414 4870
rect 2761 4378 2817 4380
rect 2841 4378 2897 4380
rect 2921 4378 2977 4380
rect 3001 4378 3057 4380
rect 2761 4326 2807 4378
rect 2807 4326 2817 4378
rect 2841 4326 2871 4378
rect 2871 4326 2883 4378
rect 2883 4326 2897 4378
rect 2921 4326 2935 4378
rect 2935 4326 2947 4378
rect 2947 4326 2977 4378
rect 3001 4326 3011 4378
rect 3011 4326 3057 4378
rect 2761 4324 2817 4326
rect 2841 4324 2897 4326
rect 2921 4324 2977 4326
rect 3001 4324 3057 4326
rect 2761 3290 2817 3292
rect 2841 3290 2897 3292
rect 2921 3290 2977 3292
rect 3001 3290 3057 3292
rect 2761 3238 2807 3290
rect 2807 3238 2817 3290
rect 2841 3238 2871 3290
rect 2871 3238 2883 3290
rect 2883 3238 2897 3290
rect 2921 3238 2935 3290
rect 2935 3238 2947 3290
rect 2947 3238 2977 3290
rect 3001 3238 3011 3290
rect 3011 3238 3057 3290
rect 2761 3236 2817 3238
rect 2841 3236 2897 3238
rect 2921 3236 2977 3238
rect 3001 3236 3057 3238
rect 2761 2202 2817 2204
rect 2841 2202 2897 2204
rect 2921 2202 2977 2204
rect 3001 2202 3057 2204
rect 2761 2150 2807 2202
rect 2807 2150 2817 2202
rect 2841 2150 2871 2202
rect 2871 2150 2883 2202
rect 2883 2150 2897 2202
rect 2921 2150 2935 2202
rect 2935 2150 2947 2202
rect 2947 2150 2977 2202
rect 3001 2150 3011 2202
rect 3011 2150 3057 2202
rect 2761 2148 2817 2150
rect 2841 2148 2897 2150
rect 2921 2148 2977 2150
rect 3001 2148 3057 2150
rect 2761 1114 2817 1116
rect 2841 1114 2897 1116
rect 2921 1114 2977 1116
rect 3001 1114 3057 1116
rect 2761 1062 2807 1114
rect 2807 1062 2817 1114
rect 2841 1062 2871 1114
rect 2871 1062 2883 1114
rect 2883 1062 2897 1114
rect 2921 1062 2935 1114
rect 2935 1062 2947 1114
rect 2947 1062 2977 1114
rect 3001 1062 3011 1114
rect 3011 1062 3057 1114
rect 2761 1060 2817 1062
rect 2841 1060 2897 1062
rect 2921 1060 2977 1062
rect 3001 1060 3057 1062
rect 5118 3834 5174 3836
rect 5198 3834 5254 3836
rect 5278 3834 5334 3836
rect 5358 3834 5414 3836
rect 5118 3782 5164 3834
rect 5164 3782 5174 3834
rect 5198 3782 5228 3834
rect 5228 3782 5240 3834
rect 5240 3782 5254 3834
rect 5278 3782 5292 3834
rect 5292 3782 5304 3834
rect 5304 3782 5334 3834
rect 5358 3782 5368 3834
rect 5368 3782 5414 3834
rect 5118 3780 5174 3782
rect 5198 3780 5254 3782
rect 5278 3780 5334 3782
rect 5358 3780 5414 3782
rect 5118 2746 5174 2748
rect 5198 2746 5254 2748
rect 5278 2746 5334 2748
rect 5358 2746 5414 2748
rect 5118 2694 5164 2746
rect 5164 2694 5174 2746
rect 5198 2694 5228 2746
rect 5228 2694 5240 2746
rect 5240 2694 5254 2746
rect 5278 2694 5292 2746
rect 5292 2694 5304 2746
rect 5304 2694 5334 2746
rect 5358 2694 5368 2746
rect 5368 2694 5414 2746
rect 5118 2692 5174 2694
rect 5198 2692 5254 2694
rect 5278 2692 5334 2694
rect 5358 2692 5414 2694
rect 5118 1658 5174 1660
rect 5198 1658 5254 1660
rect 5278 1658 5334 1660
rect 5358 1658 5414 1660
rect 5118 1606 5164 1658
rect 5164 1606 5174 1658
rect 5198 1606 5228 1658
rect 5228 1606 5240 1658
rect 5240 1606 5254 1658
rect 5278 1606 5292 1658
rect 5292 1606 5304 1658
rect 5304 1606 5334 1658
rect 5358 1606 5368 1658
rect 5368 1606 5414 1658
rect 5118 1604 5174 1606
rect 5198 1604 5254 1606
rect 5278 1604 5334 1606
rect 5358 1604 5414 1606
rect 5118 570 5174 572
rect 5198 570 5254 572
rect 5278 570 5334 572
rect 5358 570 5414 572
rect 5118 518 5164 570
rect 5164 518 5174 570
rect 5198 518 5228 570
rect 5228 518 5240 570
rect 5240 518 5254 570
rect 5278 518 5292 570
rect 5292 518 5304 570
rect 5304 518 5334 570
rect 5358 518 5368 570
rect 5368 518 5414 570
rect 5118 516 5174 518
rect 5198 516 5254 518
rect 5278 516 5334 518
rect 5358 516 5414 518
rect 7476 9818 7532 9820
rect 7556 9818 7612 9820
rect 7636 9818 7692 9820
rect 7716 9818 7772 9820
rect 7476 9766 7522 9818
rect 7522 9766 7532 9818
rect 7556 9766 7586 9818
rect 7586 9766 7598 9818
rect 7598 9766 7612 9818
rect 7636 9766 7650 9818
rect 7650 9766 7662 9818
rect 7662 9766 7692 9818
rect 7716 9766 7726 9818
rect 7726 9766 7772 9818
rect 7476 9764 7532 9766
rect 7556 9764 7612 9766
rect 7636 9764 7692 9766
rect 7716 9764 7772 9766
rect 7476 8730 7532 8732
rect 7556 8730 7612 8732
rect 7636 8730 7692 8732
rect 7716 8730 7772 8732
rect 7476 8678 7522 8730
rect 7522 8678 7532 8730
rect 7556 8678 7586 8730
rect 7586 8678 7598 8730
rect 7598 8678 7612 8730
rect 7636 8678 7650 8730
rect 7650 8678 7662 8730
rect 7662 8678 7692 8730
rect 7716 8678 7726 8730
rect 7726 8678 7772 8730
rect 7476 8676 7532 8678
rect 7556 8676 7612 8678
rect 7636 8676 7692 8678
rect 7716 8676 7772 8678
rect 7476 7642 7532 7644
rect 7556 7642 7612 7644
rect 7636 7642 7692 7644
rect 7716 7642 7772 7644
rect 7476 7590 7522 7642
rect 7522 7590 7532 7642
rect 7556 7590 7586 7642
rect 7586 7590 7598 7642
rect 7598 7590 7612 7642
rect 7636 7590 7650 7642
rect 7650 7590 7662 7642
rect 7662 7590 7692 7642
rect 7716 7590 7726 7642
rect 7726 7590 7772 7642
rect 7476 7588 7532 7590
rect 7556 7588 7612 7590
rect 7636 7588 7692 7590
rect 7716 7588 7772 7590
rect 7476 6554 7532 6556
rect 7556 6554 7612 6556
rect 7636 6554 7692 6556
rect 7716 6554 7772 6556
rect 7476 6502 7522 6554
rect 7522 6502 7532 6554
rect 7556 6502 7586 6554
rect 7586 6502 7598 6554
rect 7598 6502 7612 6554
rect 7636 6502 7650 6554
rect 7650 6502 7662 6554
rect 7662 6502 7692 6554
rect 7716 6502 7726 6554
rect 7726 6502 7772 6554
rect 7476 6500 7532 6502
rect 7556 6500 7612 6502
rect 7636 6500 7692 6502
rect 7716 6500 7772 6502
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 10073 19066 10129 19068
rect 9833 19014 9879 19066
rect 9879 19014 9889 19066
rect 9913 19014 9943 19066
rect 9943 19014 9955 19066
rect 9955 19014 9969 19066
rect 9993 19014 10007 19066
rect 10007 19014 10019 19066
rect 10019 19014 10049 19066
rect 10073 19014 10083 19066
rect 10083 19014 10129 19066
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 10073 19012 10129 19014
rect 14548 19066 14604 19068
rect 14628 19066 14684 19068
rect 14708 19066 14764 19068
rect 14788 19066 14844 19068
rect 14548 19014 14594 19066
rect 14594 19014 14604 19066
rect 14628 19014 14658 19066
rect 14658 19014 14670 19066
rect 14670 19014 14684 19066
rect 14708 19014 14722 19066
rect 14722 19014 14734 19066
rect 14734 19014 14764 19066
rect 14788 19014 14798 19066
rect 14798 19014 14844 19066
rect 14548 19012 14604 19014
rect 14628 19012 14684 19014
rect 14708 19012 14764 19014
rect 14788 19012 14844 19014
rect 8850 16632 8906 16688
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 10073 17978 10129 17980
rect 9833 17926 9879 17978
rect 9879 17926 9889 17978
rect 9913 17926 9943 17978
rect 9943 17926 9955 17978
rect 9955 17926 9969 17978
rect 9993 17926 10007 17978
rect 10007 17926 10019 17978
rect 10019 17926 10049 17978
rect 10073 17926 10083 17978
rect 10083 17926 10129 17978
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10073 17924 10129 17926
rect 12191 18522 12247 18524
rect 12271 18522 12327 18524
rect 12351 18522 12407 18524
rect 12431 18522 12487 18524
rect 12191 18470 12237 18522
rect 12237 18470 12247 18522
rect 12271 18470 12301 18522
rect 12301 18470 12313 18522
rect 12313 18470 12327 18522
rect 12351 18470 12365 18522
rect 12365 18470 12377 18522
rect 12377 18470 12407 18522
rect 12431 18470 12441 18522
rect 12441 18470 12487 18522
rect 12191 18468 12247 18470
rect 12271 18468 12327 18470
rect 12351 18468 12407 18470
rect 12431 18468 12487 18470
rect 8666 15408 8722 15464
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 10073 16890 10129 16892
rect 9833 16838 9879 16890
rect 9879 16838 9889 16890
rect 9913 16838 9943 16890
rect 9943 16838 9955 16890
rect 9955 16838 9969 16890
rect 9993 16838 10007 16890
rect 10007 16838 10019 16890
rect 10019 16838 10049 16890
rect 10073 16838 10083 16890
rect 10083 16838 10129 16890
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10073 16836 10129 16838
rect 9954 16668 9956 16688
rect 9956 16668 10008 16688
rect 10008 16668 10010 16688
rect 9954 16632 10010 16668
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 10073 15802 10129 15804
rect 9833 15750 9879 15802
rect 9879 15750 9889 15802
rect 9913 15750 9943 15802
rect 9943 15750 9955 15802
rect 9955 15750 9969 15802
rect 9993 15750 10007 15802
rect 10007 15750 10019 15802
rect 10019 15750 10049 15802
rect 10073 15750 10083 15802
rect 10083 15750 10129 15802
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 10073 15748 10129 15750
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 10073 14714 10129 14716
rect 9833 14662 9879 14714
rect 9879 14662 9889 14714
rect 9913 14662 9943 14714
rect 9943 14662 9955 14714
rect 9955 14662 9969 14714
rect 9993 14662 10007 14714
rect 10007 14662 10019 14714
rect 10019 14662 10049 14714
rect 10073 14662 10083 14714
rect 10083 14662 10129 14714
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 10073 14660 10129 14662
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 10073 13626 10129 13628
rect 9833 13574 9879 13626
rect 9879 13574 9889 13626
rect 9913 13574 9943 13626
rect 9943 13574 9955 13626
rect 9955 13574 9969 13626
rect 9993 13574 10007 13626
rect 10007 13574 10019 13626
rect 10019 13574 10049 13626
rect 10073 13574 10083 13626
rect 10083 13574 10129 13626
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10073 13572 10129 13574
rect 9586 12688 9642 12744
rect 7476 5466 7532 5468
rect 7556 5466 7612 5468
rect 7636 5466 7692 5468
rect 7716 5466 7772 5468
rect 7476 5414 7522 5466
rect 7522 5414 7532 5466
rect 7556 5414 7586 5466
rect 7586 5414 7598 5466
rect 7598 5414 7612 5466
rect 7636 5414 7650 5466
rect 7650 5414 7662 5466
rect 7662 5414 7692 5466
rect 7716 5414 7726 5466
rect 7726 5414 7772 5466
rect 7476 5412 7532 5414
rect 7556 5412 7612 5414
rect 7636 5412 7692 5414
rect 7716 5412 7772 5414
rect 7476 4378 7532 4380
rect 7556 4378 7612 4380
rect 7636 4378 7692 4380
rect 7716 4378 7772 4380
rect 7476 4326 7522 4378
rect 7522 4326 7532 4378
rect 7556 4326 7586 4378
rect 7586 4326 7598 4378
rect 7598 4326 7612 4378
rect 7636 4326 7650 4378
rect 7650 4326 7662 4378
rect 7662 4326 7692 4378
rect 7716 4326 7726 4378
rect 7726 4326 7772 4378
rect 7476 4324 7532 4326
rect 7556 4324 7612 4326
rect 7636 4324 7692 4326
rect 7716 4324 7772 4326
rect 7476 3290 7532 3292
rect 7556 3290 7612 3292
rect 7636 3290 7692 3292
rect 7716 3290 7772 3292
rect 7476 3238 7522 3290
rect 7522 3238 7532 3290
rect 7556 3238 7586 3290
rect 7586 3238 7598 3290
rect 7598 3238 7612 3290
rect 7636 3238 7650 3290
rect 7650 3238 7662 3290
rect 7662 3238 7692 3290
rect 7716 3238 7726 3290
rect 7726 3238 7772 3290
rect 7476 3236 7532 3238
rect 7556 3236 7612 3238
rect 7636 3236 7692 3238
rect 7716 3236 7772 3238
rect 7476 2202 7532 2204
rect 7556 2202 7612 2204
rect 7636 2202 7692 2204
rect 7716 2202 7772 2204
rect 7476 2150 7522 2202
rect 7522 2150 7532 2202
rect 7556 2150 7586 2202
rect 7586 2150 7598 2202
rect 7598 2150 7612 2202
rect 7636 2150 7650 2202
rect 7650 2150 7662 2202
rect 7662 2150 7692 2202
rect 7716 2150 7726 2202
rect 7726 2150 7772 2202
rect 7476 2148 7532 2150
rect 7556 2148 7612 2150
rect 7636 2148 7692 2150
rect 7716 2148 7772 2150
rect 7476 1114 7532 1116
rect 7556 1114 7612 1116
rect 7636 1114 7692 1116
rect 7716 1114 7772 1116
rect 7476 1062 7522 1114
rect 7522 1062 7532 1114
rect 7556 1062 7586 1114
rect 7586 1062 7598 1114
rect 7598 1062 7612 1114
rect 7636 1062 7650 1114
rect 7650 1062 7662 1114
rect 7662 1062 7692 1114
rect 7716 1062 7726 1114
rect 7726 1062 7772 1114
rect 7476 1060 7532 1062
rect 7556 1060 7612 1062
rect 7636 1060 7692 1062
rect 7716 1060 7772 1062
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 10073 12538 10129 12540
rect 9833 12486 9879 12538
rect 9879 12486 9889 12538
rect 9913 12486 9943 12538
rect 9943 12486 9955 12538
rect 9955 12486 9969 12538
rect 9993 12486 10007 12538
rect 10007 12486 10019 12538
rect 10019 12486 10049 12538
rect 10073 12486 10083 12538
rect 10083 12486 10129 12538
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 10073 12484 10129 12486
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 10073 11450 10129 11452
rect 9833 11398 9879 11450
rect 9879 11398 9889 11450
rect 9913 11398 9943 11450
rect 9943 11398 9955 11450
rect 9955 11398 9969 11450
rect 9993 11398 10007 11450
rect 10007 11398 10019 11450
rect 10019 11398 10049 11450
rect 10073 11398 10083 11450
rect 10083 11398 10129 11450
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 10073 11396 10129 11398
rect 10598 11736 10654 11792
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 10073 10362 10129 10364
rect 9833 10310 9879 10362
rect 9879 10310 9889 10362
rect 9913 10310 9943 10362
rect 9943 10310 9955 10362
rect 9955 10310 9969 10362
rect 9993 10310 10007 10362
rect 10007 10310 10019 10362
rect 10019 10310 10049 10362
rect 10073 10310 10083 10362
rect 10083 10310 10129 10362
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 10073 10308 10129 10310
rect 10046 9560 10102 9616
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 10073 9274 10129 9276
rect 9833 9222 9879 9274
rect 9879 9222 9889 9274
rect 9913 9222 9943 9274
rect 9943 9222 9955 9274
rect 9955 9222 9969 9274
rect 9993 9222 10007 9274
rect 10007 9222 10019 9274
rect 10019 9222 10049 9274
rect 10073 9222 10083 9274
rect 10083 9222 10129 9274
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 10073 9220 10129 9222
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 10073 8186 10129 8188
rect 9833 8134 9879 8186
rect 9879 8134 9889 8186
rect 9913 8134 9943 8186
rect 9943 8134 9955 8186
rect 9955 8134 9969 8186
rect 9993 8134 10007 8186
rect 10007 8134 10019 8186
rect 10019 8134 10049 8186
rect 10073 8134 10083 8186
rect 10083 8134 10129 8186
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 10073 8132 10129 8134
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 10073 7098 10129 7100
rect 9833 7046 9879 7098
rect 9879 7046 9889 7098
rect 9913 7046 9943 7098
rect 9943 7046 9955 7098
rect 9955 7046 9969 7098
rect 9993 7046 10007 7098
rect 10007 7046 10019 7098
rect 10019 7046 10049 7098
rect 10073 7046 10083 7098
rect 10083 7046 10129 7098
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 10073 7044 10129 7046
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 10073 6010 10129 6012
rect 9833 5958 9879 6010
rect 9879 5958 9889 6010
rect 9913 5958 9943 6010
rect 9943 5958 9955 6010
rect 9955 5958 9969 6010
rect 9993 5958 10007 6010
rect 10007 5958 10019 6010
rect 10019 5958 10049 6010
rect 10073 5958 10083 6010
rect 10083 5958 10129 6010
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10073 5956 10129 5958
rect 12191 17434 12247 17436
rect 12271 17434 12327 17436
rect 12351 17434 12407 17436
rect 12431 17434 12487 17436
rect 12191 17382 12237 17434
rect 12237 17382 12247 17434
rect 12271 17382 12301 17434
rect 12301 17382 12313 17434
rect 12313 17382 12327 17434
rect 12351 17382 12365 17434
rect 12365 17382 12377 17434
rect 12377 17382 12407 17434
rect 12431 17382 12441 17434
rect 12441 17382 12487 17434
rect 12191 17380 12247 17382
rect 12271 17380 12327 17382
rect 12351 17380 12407 17382
rect 12431 17380 12487 17382
rect 12191 16346 12247 16348
rect 12271 16346 12327 16348
rect 12351 16346 12407 16348
rect 12431 16346 12487 16348
rect 12191 16294 12237 16346
rect 12237 16294 12247 16346
rect 12271 16294 12301 16346
rect 12301 16294 12313 16346
rect 12313 16294 12327 16346
rect 12351 16294 12365 16346
rect 12365 16294 12377 16346
rect 12377 16294 12407 16346
rect 12431 16294 12441 16346
rect 12441 16294 12487 16346
rect 12191 16292 12247 16294
rect 12271 16292 12327 16294
rect 12351 16292 12407 16294
rect 12431 16292 12487 16294
rect 14548 17978 14604 17980
rect 14628 17978 14684 17980
rect 14708 17978 14764 17980
rect 14788 17978 14844 17980
rect 14548 17926 14594 17978
rect 14594 17926 14604 17978
rect 14628 17926 14658 17978
rect 14658 17926 14670 17978
rect 14670 17926 14684 17978
rect 14708 17926 14722 17978
rect 14722 17926 14734 17978
rect 14734 17926 14764 17978
rect 14788 17926 14798 17978
rect 14798 17926 14844 17978
rect 14548 17924 14604 17926
rect 14628 17924 14684 17926
rect 14708 17924 14764 17926
rect 14788 17924 14844 17926
rect 16906 18522 16962 18524
rect 16986 18522 17042 18524
rect 17066 18522 17122 18524
rect 17146 18522 17202 18524
rect 16906 18470 16952 18522
rect 16952 18470 16962 18522
rect 16986 18470 17016 18522
rect 17016 18470 17028 18522
rect 17028 18470 17042 18522
rect 17066 18470 17080 18522
rect 17080 18470 17092 18522
rect 17092 18470 17122 18522
rect 17146 18470 17156 18522
rect 17156 18470 17202 18522
rect 16906 18468 16962 18470
rect 16986 18468 17042 18470
rect 17066 18468 17122 18470
rect 17146 18468 17202 18470
rect 12191 15258 12247 15260
rect 12271 15258 12327 15260
rect 12351 15258 12407 15260
rect 12431 15258 12487 15260
rect 12191 15206 12237 15258
rect 12237 15206 12247 15258
rect 12271 15206 12301 15258
rect 12301 15206 12313 15258
rect 12313 15206 12327 15258
rect 12351 15206 12365 15258
rect 12365 15206 12377 15258
rect 12377 15206 12407 15258
rect 12431 15206 12441 15258
rect 12441 15206 12487 15258
rect 12191 15204 12247 15206
rect 12271 15204 12327 15206
rect 12351 15204 12407 15206
rect 12431 15204 12487 15206
rect 16906 17434 16962 17436
rect 16986 17434 17042 17436
rect 17066 17434 17122 17436
rect 17146 17434 17202 17436
rect 16906 17382 16952 17434
rect 16952 17382 16962 17434
rect 16986 17382 17016 17434
rect 17016 17382 17028 17434
rect 17028 17382 17042 17434
rect 17066 17382 17080 17434
rect 17080 17382 17092 17434
rect 17092 17382 17122 17434
rect 17146 17382 17156 17434
rect 17156 17382 17202 17434
rect 16906 17380 16962 17382
rect 16986 17380 17042 17382
rect 17066 17380 17122 17382
rect 17146 17380 17202 17382
rect 14548 16890 14604 16892
rect 14628 16890 14684 16892
rect 14708 16890 14764 16892
rect 14788 16890 14844 16892
rect 14548 16838 14594 16890
rect 14594 16838 14604 16890
rect 14628 16838 14658 16890
rect 14658 16838 14670 16890
rect 14670 16838 14684 16890
rect 14708 16838 14722 16890
rect 14722 16838 14734 16890
rect 14734 16838 14764 16890
rect 14788 16838 14798 16890
rect 14798 16838 14844 16890
rect 14548 16836 14604 16838
rect 14628 16836 14684 16838
rect 14708 16836 14764 16838
rect 14788 16836 14844 16838
rect 16906 16346 16962 16348
rect 16986 16346 17042 16348
rect 17066 16346 17122 16348
rect 17146 16346 17202 16348
rect 16906 16294 16952 16346
rect 16952 16294 16962 16346
rect 16986 16294 17016 16346
rect 17016 16294 17028 16346
rect 17028 16294 17042 16346
rect 17066 16294 17080 16346
rect 17080 16294 17092 16346
rect 17092 16294 17122 16346
rect 17146 16294 17156 16346
rect 17156 16294 17202 16346
rect 16906 16292 16962 16294
rect 16986 16292 17042 16294
rect 17066 16292 17122 16294
rect 17146 16292 17202 16294
rect 19263 19066 19319 19068
rect 19343 19066 19399 19068
rect 19423 19066 19479 19068
rect 19503 19066 19559 19068
rect 19263 19014 19309 19066
rect 19309 19014 19319 19066
rect 19343 19014 19373 19066
rect 19373 19014 19385 19066
rect 19385 19014 19399 19066
rect 19423 19014 19437 19066
rect 19437 19014 19449 19066
rect 19449 19014 19479 19066
rect 19503 19014 19513 19066
rect 19513 19014 19559 19066
rect 19263 19012 19319 19014
rect 19343 19012 19399 19014
rect 19423 19012 19479 19014
rect 19503 19012 19559 19014
rect 19263 17978 19319 17980
rect 19343 17978 19399 17980
rect 19423 17978 19479 17980
rect 19503 17978 19559 17980
rect 19263 17926 19309 17978
rect 19309 17926 19319 17978
rect 19343 17926 19373 17978
rect 19373 17926 19385 17978
rect 19385 17926 19399 17978
rect 19423 17926 19437 17978
rect 19437 17926 19449 17978
rect 19449 17926 19479 17978
rect 19503 17926 19513 17978
rect 19513 17926 19559 17978
rect 19263 17924 19319 17926
rect 19343 17924 19399 17926
rect 19423 17924 19479 17926
rect 19503 17924 19559 17926
rect 19263 16890 19319 16892
rect 19343 16890 19399 16892
rect 19423 16890 19479 16892
rect 19503 16890 19559 16892
rect 19263 16838 19309 16890
rect 19309 16838 19319 16890
rect 19343 16838 19373 16890
rect 19373 16838 19385 16890
rect 19385 16838 19399 16890
rect 19423 16838 19437 16890
rect 19437 16838 19449 16890
rect 19449 16838 19479 16890
rect 19503 16838 19513 16890
rect 19513 16838 19559 16890
rect 19263 16836 19319 16838
rect 19343 16836 19399 16838
rect 19423 16836 19479 16838
rect 19503 16836 19559 16838
rect 19062 15952 19118 16008
rect 14548 15802 14604 15804
rect 14628 15802 14684 15804
rect 14708 15802 14764 15804
rect 14788 15802 14844 15804
rect 14548 15750 14594 15802
rect 14594 15750 14604 15802
rect 14628 15750 14658 15802
rect 14658 15750 14670 15802
rect 14670 15750 14684 15802
rect 14708 15750 14722 15802
rect 14722 15750 14734 15802
rect 14734 15750 14764 15802
rect 14788 15750 14798 15802
rect 14798 15750 14844 15802
rect 14548 15748 14604 15750
rect 14628 15748 14684 15750
rect 14708 15748 14764 15750
rect 14788 15748 14844 15750
rect 14548 14714 14604 14716
rect 14628 14714 14684 14716
rect 14708 14714 14764 14716
rect 14788 14714 14844 14716
rect 14548 14662 14594 14714
rect 14594 14662 14604 14714
rect 14628 14662 14658 14714
rect 14658 14662 14670 14714
rect 14670 14662 14684 14714
rect 14708 14662 14722 14714
rect 14722 14662 14734 14714
rect 14734 14662 14764 14714
rect 14788 14662 14798 14714
rect 14798 14662 14844 14714
rect 14548 14660 14604 14662
rect 14628 14660 14684 14662
rect 14708 14660 14764 14662
rect 14788 14660 14844 14662
rect 19263 15802 19319 15804
rect 19343 15802 19399 15804
rect 19423 15802 19479 15804
rect 19503 15802 19559 15804
rect 19263 15750 19309 15802
rect 19309 15750 19319 15802
rect 19343 15750 19373 15802
rect 19373 15750 19385 15802
rect 19385 15750 19399 15802
rect 19423 15750 19437 15802
rect 19437 15750 19449 15802
rect 19449 15750 19479 15802
rect 19503 15750 19513 15802
rect 19513 15750 19559 15802
rect 19263 15748 19319 15750
rect 19343 15748 19399 15750
rect 19423 15748 19479 15750
rect 19503 15748 19559 15750
rect 16906 15258 16962 15260
rect 16986 15258 17042 15260
rect 17066 15258 17122 15260
rect 17146 15258 17202 15260
rect 16906 15206 16952 15258
rect 16952 15206 16962 15258
rect 16986 15206 17016 15258
rect 17016 15206 17028 15258
rect 17028 15206 17042 15258
rect 17066 15206 17080 15258
rect 17080 15206 17092 15258
rect 17092 15206 17122 15258
rect 17146 15206 17156 15258
rect 17156 15206 17202 15258
rect 16906 15204 16962 15206
rect 16986 15204 17042 15206
rect 17066 15204 17122 15206
rect 17146 15204 17202 15206
rect 12191 14170 12247 14172
rect 12271 14170 12327 14172
rect 12351 14170 12407 14172
rect 12431 14170 12487 14172
rect 12191 14118 12237 14170
rect 12237 14118 12247 14170
rect 12271 14118 12301 14170
rect 12301 14118 12313 14170
rect 12313 14118 12327 14170
rect 12351 14118 12365 14170
rect 12365 14118 12377 14170
rect 12377 14118 12407 14170
rect 12431 14118 12441 14170
rect 12441 14118 12487 14170
rect 12191 14116 12247 14118
rect 12271 14116 12327 14118
rect 12351 14116 12407 14118
rect 12431 14116 12487 14118
rect 12191 13082 12247 13084
rect 12271 13082 12327 13084
rect 12351 13082 12407 13084
rect 12431 13082 12487 13084
rect 12191 13030 12237 13082
rect 12237 13030 12247 13082
rect 12271 13030 12301 13082
rect 12301 13030 12313 13082
rect 12313 13030 12327 13082
rect 12351 13030 12365 13082
rect 12365 13030 12377 13082
rect 12377 13030 12407 13082
rect 12431 13030 12441 13082
rect 12441 13030 12487 13082
rect 12191 13028 12247 13030
rect 12271 13028 12327 13030
rect 12351 13028 12407 13030
rect 12431 13028 12487 13030
rect 11518 12708 11574 12744
rect 11518 12688 11520 12708
rect 11520 12688 11572 12708
rect 11572 12688 11574 12708
rect 14548 13626 14604 13628
rect 14628 13626 14684 13628
rect 14708 13626 14764 13628
rect 14788 13626 14844 13628
rect 14548 13574 14594 13626
rect 14594 13574 14604 13626
rect 14628 13574 14658 13626
rect 14658 13574 14670 13626
rect 14670 13574 14684 13626
rect 14708 13574 14722 13626
rect 14722 13574 14734 13626
rect 14734 13574 14764 13626
rect 14788 13574 14798 13626
rect 14798 13574 14844 13626
rect 14548 13572 14604 13574
rect 14628 13572 14684 13574
rect 14708 13572 14764 13574
rect 14788 13572 14844 13574
rect 14548 12538 14604 12540
rect 14628 12538 14684 12540
rect 14708 12538 14764 12540
rect 14788 12538 14844 12540
rect 14548 12486 14594 12538
rect 14594 12486 14604 12538
rect 14628 12486 14658 12538
rect 14658 12486 14670 12538
rect 14670 12486 14684 12538
rect 14708 12486 14722 12538
rect 14722 12486 14734 12538
rect 14734 12486 14764 12538
rect 14788 12486 14798 12538
rect 14798 12486 14844 12538
rect 14548 12484 14604 12486
rect 14628 12484 14684 12486
rect 14708 12484 14764 12486
rect 14788 12484 14844 12486
rect 12191 11994 12247 11996
rect 12271 11994 12327 11996
rect 12351 11994 12407 11996
rect 12431 11994 12487 11996
rect 12191 11942 12237 11994
rect 12237 11942 12247 11994
rect 12271 11942 12301 11994
rect 12301 11942 12313 11994
rect 12313 11942 12327 11994
rect 12351 11942 12365 11994
rect 12365 11942 12377 11994
rect 12377 11942 12407 11994
rect 12431 11942 12441 11994
rect 12441 11942 12487 11994
rect 12191 11940 12247 11942
rect 12271 11940 12327 11942
rect 12351 11940 12407 11942
rect 12431 11940 12487 11942
rect 12191 10906 12247 10908
rect 12271 10906 12327 10908
rect 12351 10906 12407 10908
rect 12431 10906 12487 10908
rect 12191 10854 12237 10906
rect 12237 10854 12247 10906
rect 12271 10854 12301 10906
rect 12301 10854 12313 10906
rect 12313 10854 12327 10906
rect 12351 10854 12365 10906
rect 12365 10854 12377 10906
rect 12377 10854 12407 10906
rect 12431 10854 12441 10906
rect 12441 10854 12487 10906
rect 12191 10852 12247 10854
rect 12271 10852 12327 10854
rect 12351 10852 12407 10854
rect 12431 10852 12487 10854
rect 10782 9560 10838 9616
rect 12191 9818 12247 9820
rect 12271 9818 12327 9820
rect 12351 9818 12407 9820
rect 12431 9818 12487 9820
rect 12191 9766 12237 9818
rect 12237 9766 12247 9818
rect 12271 9766 12301 9818
rect 12301 9766 12313 9818
rect 12313 9766 12327 9818
rect 12351 9766 12365 9818
rect 12365 9766 12377 9818
rect 12377 9766 12407 9818
rect 12431 9766 12441 9818
rect 12441 9766 12487 9818
rect 12191 9764 12247 9766
rect 12271 9764 12327 9766
rect 12351 9764 12407 9766
rect 12431 9764 12487 9766
rect 12191 8730 12247 8732
rect 12271 8730 12327 8732
rect 12351 8730 12407 8732
rect 12431 8730 12487 8732
rect 12191 8678 12237 8730
rect 12237 8678 12247 8730
rect 12271 8678 12301 8730
rect 12301 8678 12313 8730
rect 12313 8678 12327 8730
rect 12351 8678 12365 8730
rect 12365 8678 12377 8730
rect 12377 8678 12407 8730
rect 12431 8678 12441 8730
rect 12441 8678 12487 8730
rect 12191 8676 12247 8678
rect 12271 8676 12327 8678
rect 12351 8676 12407 8678
rect 12431 8676 12487 8678
rect 13082 10104 13138 10160
rect 12191 7642 12247 7644
rect 12271 7642 12327 7644
rect 12351 7642 12407 7644
rect 12431 7642 12487 7644
rect 12191 7590 12237 7642
rect 12237 7590 12247 7642
rect 12271 7590 12301 7642
rect 12301 7590 12313 7642
rect 12313 7590 12327 7642
rect 12351 7590 12365 7642
rect 12365 7590 12377 7642
rect 12377 7590 12407 7642
rect 12431 7590 12441 7642
rect 12441 7590 12487 7642
rect 12191 7588 12247 7590
rect 12271 7588 12327 7590
rect 12351 7588 12407 7590
rect 12431 7588 12487 7590
rect 11150 6860 11206 6896
rect 11150 6840 11152 6860
rect 11152 6840 11204 6860
rect 11204 6840 11206 6860
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 10073 4922 10129 4924
rect 9833 4870 9879 4922
rect 9879 4870 9889 4922
rect 9913 4870 9943 4922
rect 9943 4870 9955 4922
rect 9955 4870 9969 4922
rect 9993 4870 10007 4922
rect 10007 4870 10019 4922
rect 10019 4870 10049 4922
rect 10073 4870 10083 4922
rect 10083 4870 10129 4922
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 10073 4868 10129 4870
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 10073 3834 10129 3836
rect 9833 3782 9879 3834
rect 9879 3782 9889 3834
rect 9913 3782 9943 3834
rect 9943 3782 9955 3834
rect 9955 3782 9969 3834
rect 9993 3782 10007 3834
rect 10007 3782 10019 3834
rect 10019 3782 10049 3834
rect 10073 3782 10083 3834
rect 10083 3782 10129 3834
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 10073 3780 10129 3782
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 10073 2746 10129 2748
rect 9833 2694 9879 2746
rect 9879 2694 9889 2746
rect 9913 2694 9943 2746
rect 9943 2694 9955 2746
rect 9955 2694 9969 2746
rect 9993 2694 10007 2746
rect 10007 2694 10019 2746
rect 10019 2694 10049 2746
rect 10073 2694 10083 2746
rect 10083 2694 10129 2746
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10073 2692 10129 2694
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 10073 1658 10129 1660
rect 9833 1606 9879 1658
rect 9879 1606 9889 1658
rect 9913 1606 9943 1658
rect 9943 1606 9955 1658
rect 9955 1606 9969 1658
rect 9993 1606 10007 1658
rect 10007 1606 10019 1658
rect 10019 1606 10049 1658
rect 10073 1606 10083 1658
rect 10083 1606 10129 1658
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 10073 1604 10129 1606
rect 9833 570 9889 572
rect 9913 570 9969 572
rect 9993 570 10049 572
rect 10073 570 10129 572
rect 9833 518 9879 570
rect 9879 518 9889 570
rect 9913 518 9943 570
rect 9943 518 9955 570
rect 9955 518 9969 570
rect 9993 518 10007 570
rect 10007 518 10019 570
rect 10019 518 10049 570
rect 10073 518 10083 570
rect 10083 518 10129 570
rect 9833 516 9889 518
rect 9913 516 9969 518
rect 9993 516 10049 518
rect 10073 516 10129 518
rect 13634 10260 13690 10296
rect 13634 10240 13636 10260
rect 13636 10240 13688 10260
rect 13688 10240 13690 10260
rect 13634 9968 13690 10024
rect 14548 11450 14604 11452
rect 14628 11450 14684 11452
rect 14708 11450 14764 11452
rect 14788 11450 14844 11452
rect 14548 11398 14594 11450
rect 14594 11398 14604 11450
rect 14628 11398 14658 11450
rect 14658 11398 14670 11450
rect 14670 11398 14684 11450
rect 14708 11398 14722 11450
rect 14722 11398 14734 11450
rect 14734 11398 14764 11450
rect 14788 11398 14798 11450
rect 14798 11398 14844 11450
rect 14548 11396 14604 11398
rect 14628 11396 14684 11398
rect 14708 11396 14764 11398
rect 14788 11396 14844 11398
rect 14548 10362 14604 10364
rect 14628 10362 14684 10364
rect 14708 10362 14764 10364
rect 14788 10362 14844 10364
rect 14548 10310 14594 10362
rect 14594 10310 14604 10362
rect 14628 10310 14658 10362
rect 14658 10310 14670 10362
rect 14670 10310 14684 10362
rect 14708 10310 14722 10362
rect 14722 10310 14734 10362
rect 14734 10310 14764 10362
rect 14788 10310 14798 10362
rect 14798 10310 14844 10362
rect 14548 10308 14604 10310
rect 14628 10308 14684 10310
rect 14708 10308 14764 10310
rect 14788 10308 14844 10310
rect 14370 10240 14426 10296
rect 14186 10104 14242 10160
rect 14738 9988 14794 10024
rect 14738 9968 14740 9988
rect 14740 9968 14792 9988
rect 14792 9968 14794 9988
rect 14548 9274 14604 9276
rect 14628 9274 14684 9276
rect 14708 9274 14764 9276
rect 14788 9274 14844 9276
rect 14548 9222 14594 9274
rect 14594 9222 14604 9274
rect 14628 9222 14658 9274
rect 14658 9222 14670 9274
rect 14670 9222 14684 9274
rect 14708 9222 14722 9274
rect 14722 9222 14734 9274
rect 14734 9222 14764 9274
rect 14788 9222 14798 9274
rect 14798 9222 14844 9274
rect 14548 9220 14604 9222
rect 14628 9220 14684 9222
rect 14708 9220 14764 9222
rect 14788 9220 14844 9222
rect 19263 14714 19319 14716
rect 19343 14714 19399 14716
rect 19423 14714 19479 14716
rect 19503 14714 19559 14716
rect 19263 14662 19309 14714
rect 19309 14662 19319 14714
rect 19343 14662 19373 14714
rect 19373 14662 19385 14714
rect 19385 14662 19399 14714
rect 19423 14662 19437 14714
rect 19437 14662 19449 14714
rect 19449 14662 19479 14714
rect 19503 14662 19513 14714
rect 19513 14662 19559 14714
rect 19263 14660 19319 14662
rect 19343 14660 19399 14662
rect 19423 14660 19479 14662
rect 19503 14660 19559 14662
rect 16906 14170 16962 14172
rect 16986 14170 17042 14172
rect 17066 14170 17122 14172
rect 17146 14170 17202 14172
rect 16906 14118 16952 14170
rect 16952 14118 16962 14170
rect 16986 14118 17016 14170
rect 17016 14118 17028 14170
rect 17028 14118 17042 14170
rect 17066 14118 17080 14170
rect 17080 14118 17092 14170
rect 17092 14118 17122 14170
rect 17146 14118 17156 14170
rect 17156 14118 17202 14170
rect 16906 14116 16962 14118
rect 16986 14116 17042 14118
rect 17066 14116 17122 14118
rect 17146 14116 17202 14118
rect 19263 13626 19319 13628
rect 19343 13626 19399 13628
rect 19423 13626 19479 13628
rect 19503 13626 19559 13628
rect 19263 13574 19309 13626
rect 19309 13574 19319 13626
rect 19343 13574 19373 13626
rect 19373 13574 19385 13626
rect 19385 13574 19399 13626
rect 19423 13574 19437 13626
rect 19437 13574 19449 13626
rect 19449 13574 19479 13626
rect 19503 13574 19513 13626
rect 19513 13574 19559 13626
rect 19263 13572 19319 13574
rect 19343 13572 19399 13574
rect 19423 13572 19479 13574
rect 19503 13572 19559 13574
rect 16906 13082 16962 13084
rect 16986 13082 17042 13084
rect 17066 13082 17122 13084
rect 17146 13082 17202 13084
rect 16906 13030 16952 13082
rect 16952 13030 16962 13082
rect 16986 13030 17016 13082
rect 17016 13030 17028 13082
rect 17028 13030 17042 13082
rect 17066 13030 17080 13082
rect 17080 13030 17092 13082
rect 17092 13030 17122 13082
rect 17146 13030 17156 13082
rect 17156 13030 17202 13082
rect 16906 13028 16962 13030
rect 16986 13028 17042 13030
rect 17066 13028 17122 13030
rect 17146 13028 17202 13030
rect 16906 11994 16962 11996
rect 16986 11994 17042 11996
rect 17066 11994 17122 11996
rect 17146 11994 17202 11996
rect 16906 11942 16952 11994
rect 16952 11942 16962 11994
rect 16986 11942 17016 11994
rect 17016 11942 17028 11994
rect 17028 11942 17042 11994
rect 17066 11942 17080 11994
rect 17080 11942 17092 11994
rect 17092 11942 17122 11994
rect 17146 11942 17156 11994
rect 17156 11942 17202 11994
rect 16906 11940 16962 11942
rect 16986 11940 17042 11942
rect 17066 11940 17122 11942
rect 17146 11940 17202 11942
rect 14548 8186 14604 8188
rect 14628 8186 14684 8188
rect 14708 8186 14764 8188
rect 14788 8186 14844 8188
rect 14548 8134 14594 8186
rect 14594 8134 14604 8186
rect 14628 8134 14658 8186
rect 14658 8134 14670 8186
rect 14670 8134 14684 8186
rect 14708 8134 14722 8186
rect 14722 8134 14734 8186
rect 14734 8134 14764 8186
rect 14788 8134 14798 8186
rect 14798 8134 14844 8186
rect 14548 8132 14604 8134
rect 14628 8132 14684 8134
rect 14708 8132 14764 8134
rect 14788 8132 14844 8134
rect 14548 7098 14604 7100
rect 14628 7098 14684 7100
rect 14708 7098 14764 7100
rect 14788 7098 14844 7100
rect 14548 7046 14594 7098
rect 14594 7046 14604 7098
rect 14628 7046 14658 7098
rect 14658 7046 14670 7098
rect 14670 7046 14684 7098
rect 14708 7046 14722 7098
rect 14722 7046 14734 7098
rect 14734 7046 14764 7098
rect 14788 7046 14798 7098
rect 14798 7046 14844 7098
rect 14548 7044 14604 7046
rect 14628 7044 14684 7046
rect 14708 7044 14764 7046
rect 14788 7044 14844 7046
rect 16906 10906 16962 10908
rect 16986 10906 17042 10908
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 16906 10854 16952 10906
rect 16952 10854 16962 10906
rect 16986 10854 17016 10906
rect 17016 10854 17028 10906
rect 17028 10854 17042 10906
rect 17066 10854 17080 10906
rect 17080 10854 17092 10906
rect 17092 10854 17122 10906
rect 17146 10854 17156 10906
rect 17156 10854 17202 10906
rect 16906 10852 16962 10854
rect 16986 10852 17042 10854
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 12191 6554 12247 6556
rect 12271 6554 12327 6556
rect 12351 6554 12407 6556
rect 12431 6554 12487 6556
rect 12191 6502 12237 6554
rect 12237 6502 12247 6554
rect 12271 6502 12301 6554
rect 12301 6502 12313 6554
rect 12313 6502 12327 6554
rect 12351 6502 12365 6554
rect 12365 6502 12377 6554
rect 12377 6502 12407 6554
rect 12431 6502 12441 6554
rect 12441 6502 12487 6554
rect 12191 6500 12247 6502
rect 12271 6500 12327 6502
rect 12351 6500 12407 6502
rect 12431 6500 12487 6502
rect 16906 9818 16962 9820
rect 16986 9818 17042 9820
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 16906 9766 16952 9818
rect 16952 9766 16962 9818
rect 16986 9766 17016 9818
rect 17016 9766 17028 9818
rect 17028 9766 17042 9818
rect 17066 9766 17080 9818
rect 17080 9766 17092 9818
rect 17092 9766 17122 9818
rect 17146 9766 17156 9818
rect 17156 9766 17202 9818
rect 16906 9764 16962 9766
rect 16986 9764 17042 9766
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 16906 8730 16962 8732
rect 16986 8730 17042 8732
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 16906 8678 16952 8730
rect 16952 8678 16962 8730
rect 16986 8678 17016 8730
rect 17016 8678 17028 8730
rect 17028 8678 17042 8730
rect 17066 8678 17080 8730
rect 17080 8678 17092 8730
rect 17092 8678 17122 8730
rect 17146 8678 17156 8730
rect 17156 8678 17202 8730
rect 16906 8676 16962 8678
rect 16986 8676 17042 8678
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 14548 6010 14604 6012
rect 14628 6010 14684 6012
rect 14708 6010 14764 6012
rect 14788 6010 14844 6012
rect 14548 5958 14594 6010
rect 14594 5958 14604 6010
rect 14628 5958 14658 6010
rect 14658 5958 14670 6010
rect 14670 5958 14684 6010
rect 14708 5958 14722 6010
rect 14722 5958 14734 6010
rect 14734 5958 14764 6010
rect 14788 5958 14798 6010
rect 14798 5958 14844 6010
rect 14548 5956 14604 5958
rect 14628 5956 14684 5958
rect 14708 5956 14764 5958
rect 14788 5956 14844 5958
rect 16906 7642 16962 7644
rect 16986 7642 17042 7644
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 16906 7590 16952 7642
rect 16952 7590 16962 7642
rect 16986 7590 17016 7642
rect 17016 7590 17028 7642
rect 17028 7590 17042 7642
rect 17066 7590 17080 7642
rect 17080 7590 17092 7642
rect 17092 7590 17122 7642
rect 17146 7590 17156 7642
rect 17156 7590 17202 7642
rect 16906 7588 16962 7590
rect 16986 7588 17042 7590
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 19263 12538 19319 12540
rect 19343 12538 19399 12540
rect 19423 12538 19479 12540
rect 19503 12538 19559 12540
rect 19263 12486 19309 12538
rect 19309 12486 19319 12538
rect 19343 12486 19373 12538
rect 19373 12486 19385 12538
rect 19385 12486 19399 12538
rect 19423 12486 19437 12538
rect 19437 12486 19449 12538
rect 19449 12486 19479 12538
rect 19503 12486 19513 12538
rect 19513 12486 19559 12538
rect 19263 12484 19319 12486
rect 19343 12484 19399 12486
rect 19423 12484 19479 12486
rect 19503 12484 19559 12486
rect 19263 11450 19319 11452
rect 19343 11450 19399 11452
rect 19423 11450 19479 11452
rect 19503 11450 19559 11452
rect 19263 11398 19309 11450
rect 19309 11398 19319 11450
rect 19343 11398 19373 11450
rect 19373 11398 19385 11450
rect 19385 11398 19399 11450
rect 19423 11398 19437 11450
rect 19437 11398 19449 11450
rect 19449 11398 19479 11450
rect 19503 11398 19513 11450
rect 19513 11398 19559 11450
rect 19263 11396 19319 11398
rect 19343 11396 19399 11398
rect 19423 11396 19479 11398
rect 19503 11396 19559 11398
rect 19263 10362 19319 10364
rect 19343 10362 19399 10364
rect 19423 10362 19479 10364
rect 19503 10362 19559 10364
rect 19263 10310 19309 10362
rect 19309 10310 19319 10362
rect 19343 10310 19373 10362
rect 19373 10310 19385 10362
rect 19385 10310 19399 10362
rect 19423 10310 19437 10362
rect 19437 10310 19449 10362
rect 19449 10310 19479 10362
rect 19503 10310 19513 10362
rect 19513 10310 19559 10362
rect 19263 10308 19319 10310
rect 19343 10308 19399 10310
rect 19423 10308 19479 10310
rect 19503 10308 19559 10310
rect 19263 9274 19319 9276
rect 19343 9274 19399 9276
rect 19423 9274 19479 9276
rect 19503 9274 19559 9276
rect 19263 9222 19309 9274
rect 19309 9222 19319 9274
rect 19343 9222 19373 9274
rect 19373 9222 19385 9274
rect 19385 9222 19399 9274
rect 19423 9222 19437 9274
rect 19437 9222 19449 9274
rect 19449 9222 19479 9274
rect 19503 9222 19513 9274
rect 19513 9222 19559 9274
rect 19263 9220 19319 9222
rect 19343 9220 19399 9222
rect 19423 9220 19479 9222
rect 19503 9220 19559 9222
rect 19263 8186 19319 8188
rect 19343 8186 19399 8188
rect 19423 8186 19479 8188
rect 19503 8186 19559 8188
rect 19263 8134 19309 8186
rect 19309 8134 19319 8186
rect 19343 8134 19373 8186
rect 19373 8134 19385 8186
rect 19385 8134 19399 8186
rect 19423 8134 19437 8186
rect 19437 8134 19449 8186
rect 19449 8134 19479 8186
rect 19503 8134 19513 8186
rect 19513 8134 19559 8186
rect 19263 8132 19319 8134
rect 19343 8132 19399 8134
rect 19423 8132 19479 8134
rect 19503 8132 19559 8134
rect 19263 7098 19319 7100
rect 19343 7098 19399 7100
rect 19423 7098 19479 7100
rect 19503 7098 19559 7100
rect 19263 7046 19309 7098
rect 19309 7046 19319 7098
rect 19343 7046 19373 7098
rect 19373 7046 19385 7098
rect 19385 7046 19399 7098
rect 19423 7046 19437 7098
rect 19437 7046 19449 7098
rect 19449 7046 19479 7098
rect 19503 7046 19513 7098
rect 19513 7046 19559 7098
rect 19263 7044 19319 7046
rect 19343 7044 19399 7046
rect 19423 7044 19479 7046
rect 19503 7044 19559 7046
rect 16906 6554 16962 6556
rect 16986 6554 17042 6556
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 16906 6502 16952 6554
rect 16952 6502 16962 6554
rect 16986 6502 17016 6554
rect 17016 6502 17028 6554
rect 17028 6502 17042 6554
rect 17066 6502 17080 6554
rect 17080 6502 17092 6554
rect 17092 6502 17122 6554
rect 17146 6502 17156 6554
rect 17156 6502 17202 6554
rect 16906 6500 16962 6502
rect 16986 6500 17042 6502
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 19263 6010 19319 6012
rect 19343 6010 19399 6012
rect 19423 6010 19479 6012
rect 19503 6010 19559 6012
rect 19263 5958 19309 6010
rect 19309 5958 19319 6010
rect 19343 5958 19373 6010
rect 19373 5958 19385 6010
rect 19385 5958 19399 6010
rect 19423 5958 19437 6010
rect 19437 5958 19449 6010
rect 19449 5958 19479 6010
rect 19503 5958 19513 6010
rect 19513 5958 19559 6010
rect 19263 5956 19319 5958
rect 19343 5956 19399 5958
rect 19423 5956 19479 5958
rect 19503 5956 19559 5958
rect 12191 5466 12247 5468
rect 12271 5466 12327 5468
rect 12351 5466 12407 5468
rect 12431 5466 12487 5468
rect 12191 5414 12237 5466
rect 12237 5414 12247 5466
rect 12271 5414 12301 5466
rect 12301 5414 12313 5466
rect 12313 5414 12327 5466
rect 12351 5414 12365 5466
rect 12365 5414 12377 5466
rect 12377 5414 12407 5466
rect 12431 5414 12441 5466
rect 12441 5414 12487 5466
rect 12191 5412 12247 5414
rect 12271 5412 12327 5414
rect 12351 5412 12407 5414
rect 12431 5412 12487 5414
rect 12191 4378 12247 4380
rect 12271 4378 12327 4380
rect 12351 4378 12407 4380
rect 12431 4378 12487 4380
rect 12191 4326 12237 4378
rect 12237 4326 12247 4378
rect 12271 4326 12301 4378
rect 12301 4326 12313 4378
rect 12313 4326 12327 4378
rect 12351 4326 12365 4378
rect 12365 4326 12377 4378
rect 12377 4326 12407 4378
rect 12431 4326 12441 4378
rect 12441 4326 12487 4378
rect 12191 4324 12247 4326
rect 12271 4324 12327 4326
rect 12351 4324 12407 4326
rect 12431 4324 12487 4326
rect 12191 3290 12247 3292
rect 12271 3290 12327 3292
rect 12351 3290 12407 3292
rect 12431 3290 12487 3292
rect 12191 3238 12237 3290
rect 12237 3238 12247 3290
rect 12271 3238 12301 3290
rect 12301 3238 12313 3290
rect 12313 3238 12327 3290
rect 12351 3238 12365 3290
rect 12365 3238 12377 3290
rect 12377 3238 12407 3290
rect 12431 3238 12441 3290
rect 12441 3238 12487 3290
rect 12191 3236 12247 3238
rect 12271 3236 12327 3238
rect 12351 3236 12407 3238
rect 12431 3236 12487 3238
rect 12191 2202 12247 2204
rect 12271 2202 12327 2204
rect 12351 2202 12407 2204
rect 12431 2202 12487 2204
rect 12191 2150 12237 2202
rect 12237 2150 12247 2202
rect 12271 2150 12301 2202
rect 12301 2150 12313 2202
rect 12313 2150 12327 2202
rect 12351 2150 12365 2202
rect 12365 2150 12377 2202
rect 12377 2150 12407 2202
rect 12431 2150 12441 2202
rect 12441 2150 12487 2202
rect 12191 2148 12247 2150
rect 12271 2148 12327 2150
rect 12351 2148 12407 2150
rect 12431 2148 12487 2150
rect 12191 1114 12247 1116
rect 12271 1114 12327 1116
rect 12351 1114 12407 1116
rect 12431 1114 12487 1116
rect 12191 1062 12237 1114
rect 12237 1062 12247 1114
rect 12271 1062 12301 1114
rect 12301 1062 12313 1114
rect 12313 1062 12327 1114
rect 12351 1062 12365 1114
rect 12365 1062 12377 1114
rect 12377 1062 12407 1114
rect 12431 1062 12441 1114
rect 12441 1062 12487 1114
rect 12191 1060 12247 1062
rect 12271 1060 12327 1062
rect 12351 1060 12407 1062
rect 12431 1060 12487 1062
rect 14548 4922 14604 4924
rect 14628 4922 14684 4924
rect 14708 4922 14764 4924
rect 14788 4922 14844 4924
rect 14548 4870 14594 4922
rect 14594 4870 14604 4922
rect 14628 4870 14658 4922
rect 14658 4870 14670 4922
rect 14670 4870 14684 4922
rect 14708 4870 14722 4922
rect 14722 4870 14734 4922
rect 14734 4870 14764 4922
rect 14788 4870 14798 4922
rect 14798 4870 14844 4922
rect 14548 4868 14604 4870
rect 14628 4868 14684 4870
rect 14708 4868 14764 4870
rect 14788 4868 14844 4870
rect 14548 3834 14604 3836
rect 14628 3834 14684 3836
rect 14708 3834 14764 3836
rect 14788 3834 14844 3836
rect 14548 3782 14594 3834
rect 14594 3782 14604 3834
rect 14628 3782 14658 3834
rect 14658 3782 14670 3834
rect 14670 3782 14684 3834
rect 14708 3782 14722 3834
rect 14722 3782 14734 3834
rect 14734 3782 14764 3834
rect 14788 3782 14798 3834
rect 14798 3782 14844 3834
rect 14548 3780 14604 3782
rect 14628 3780 14684 3782
rect 14708 3780 14764 3782
rect 14788 3780 14844 3782
rect 14548 2746 14604 2748
rect 14628 2746 14684 2748
rect 14708 2746 14764 2748
rect 14788 2746 14844 2748
rect 14548 2694 14594 2746
rect 14594 2694 14604 2746
rect 14628 2694 14658 2746
rect 14658 2694 14670 2746
rect 14670 2694 14684 2746
rect 14708 2694 14722 2746
rect 14722 2694 14734 2746
rect 14734 2694 14764 2746
rect 14788 2694 14798 2746
rect 14798 2694 14844 2746
rect 14548 2692 14604 2694
rect 14628 2692 14684 2694
rect 14708 2692 14764 2694
rect 14788 2692 14844 2694
rect 14548 1658 14604 1660
rect 14628 1658 14684 1660
rect 14708 1658 14764 1660
rect 14788 1658 14844 1660
rect 14548 1606 14594 1658
rect 14594 1606 14604 1658
rect 14628 1606 14658 1658
rect 14658 1606 14670 1658
rect 14670 1606 14684 1658
rect 14708 1606 14722 1658
rect 14722 1606 14734 1658
rect 14734 1606 14764 1658
rect 14788 1606 14798 1658
rect 14798 1606 14844 1658
rect 14548 1604 14604 1606
rect 14628 1604 14684 1606
rect 14708 1604 14764 1606
rect 14788 1604 14844 1606
rect 14548 570 14604 572
rect 14628 570 14684 572
rect 14708 570 14764 572
rect 14788 570 14844 572
rect 14548 518 14594 570
rect 14594 518 14604 570
rect 14628 518 14658 570
rect 14658 518 14670 570
rect 14670 518 14684 570
rect 14708 518 14722 570
rect 14722 518 14734 570
rect 14734 518 14764 570
rect 14788 518 14798 570
rect 14798 518 14844 570
rect 14548 516 14604 518
rect 14628 516 14684 518
rect 14708 516 14764 518
rect 14788 516 14844 518
rect 16906 5466 16962 5468
rect 16986 5466 17042 5468
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 16906 5414 16952 5466
rect 16952 5414 16962 5466
rect 16986 5414 17016 5466
rect 17016 5414 17028 5466
rect 17028 5414 17042 5466
rect 17066 5414 17080 5466
rect 17080 5414 17092 5466
rect 17092 5414 17122 5466
rect 17146 5414 17156 5466
rect 17156 5414 17202 5466
rect 16906 5412 16962 5414
rect 16986 5412 17042 5414
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 16906 4378 16962 4380
rect 16986 4378 17042 4380
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 16906 4326 16952 4378
rect 16952 4326 16962 4378
rect 16986 4326 17016 4378
rect 17016 4326 17028 4378
rect 17028 4326 17042 4378
rect 17066 4326 17080 4378
rect 17080 4326 17092 4378
rect 17092 4326 17122 4378
rect 17146 4326 17156 4378
rect 17156 4326 17202 4378
rect 16906 4324 16962 4326
rect 16986 4324 17042 4326
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 16906 3290 16962 3292
rect 16986 3290 17042 3292
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 16906 3238 16952 3290
rect 16952 3238 16962 3290
rect 16986 3238 17016 3290
rect 17016 3238 17028 3290
rect 17028 3238 17042 3290
rect 17066 3238 17080 3290
rect 17080 3238 17092 3290
rect 17092 3238 17122 3290
rect 17146 3238 17156 3290
rect 17156 3238 17202 3290
rect 16906 3236 16962 3238
rect 16986 3236 17042 3238
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 16906 2202 16962 2204
rect 16986 2202 17042 2204
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 16906 2150 16952 2202
rect 16952 2150 16962 2202
rect 16986 2150 17016 2202
rect 17016 2150 17028 2202
rect 17028 2150 17042 2202
rect 17066 2150 17080 2202
rect 17080 2150 17092 2202
rect 17092 2150 17122 2202
rect 17146 2150 17156 2202
rect 17156 2150 17202 2202
rect 16906 2148 16962 2150
rect 16986 2148 17042 2150
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 16906 1114 16962 1116
rect 16986 1114 17042 1116
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 16906 1062 16952 1114
rect 16952 1062 16962 1114
rect 16986 1062 17016 1114
rect 17016 1062 17028 1114
rect 17028 1062 17042 1114
rect 17066 1062 17080 1114
rect 17080 1062 17092 1114
rect 17092 1062 17122 1114
rect 17146 1062 17156 1114
rect 17156 1062 17202 1114
rect 16906 1060 16962 1062
rect 16986 1060 17042 1062
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 19263 4922 19319 4924
rect 19343 4922 19399 4924
rect 19423 4922 19479 4924
rect 19503 4922 19559 4924
rect 19263 4870 19309 4922
rect 19309 4870 19319 4922
rect 19343 4870 19373 4922
rect 19373 4870 19385 4922
rect 19385 4870 19399 4922
rect 19423 4870 19437 4922
rect 19437 4870 19449 4922
rect 19449 4870 19479 4922
rect 19503 4870 19513 4922
rect 19513 4870 19559 4922
rect 19263 4868 19319 4870
rect 19343 4868 19399 4870
rect 19423 4868 19479 4870
rect 19503 4868 19559 4870
rect 19263 3834 19319 3836
rect 19343 3834 19399 3836
rect 19423 3834 19479 3836
rect 19503 3834 19559 3836
rect 19263 3782 19309 3834
rect 19309 3782 19319 3834
rect 19343 3782 19373 3834
rect 19373 3782 19385 3834
rect 19385 3782 19399 3834
rect 19423 3782 19437 3834
rect 19437 3782 19449 3834
rect 19449 3782 19479 3834
rect 19503 3782 19513 3834
rect 19513 3782 19559 3834
rect 19263 3780 19319 3782
rect 19343 3780 19399 3782
rect 19423 3780 19479 3782
rect 19503 3780 19559 3782
rect 19263 2746 19319 2748
rect 19343 2746 19399 2748
rect 19423 2746 19479 2748
rect 19503 2746 19559 2748
rect 19263 2694 19309 2746
rect 19309 2694 19319 2746
rect 19343 2694 19373 2746
rect 19373 2694 19385 2746
rect 19385 2694 19399 2746
rect 19423 2694 19437 2746
rect 19437 2694 19449 2746
rect 19449 2694 19479 2746
rect 19503 2694 19513 2746
rect 19513 2694 19559 2746
rect 19263 2692 19319 2694
rect 19343 2692 19399 2694
rect 19423 2692 19479 2694
rect 19503 2692 19559 2694
rect 19263 1658 19319 1660
rect 19343 1658 19399 1660
rect 19423 1658 19479 1660
rect 19503 1658 19559 1660
rect 19263 1606 19309 1658
rect 19309 1606 19319 1658
rect 19343 1606 19373 1658
rect 19373 1606 19385 1658
rect 19385 1606 19399 1658
rect 19423 1606 19437 1658
rect 19437 1606 19449 1658
rect 19449 1606 19479 1658
rect 19503 1606 19513 1658
rect 19513 1606 19559 1658
rect 19263 1604 19319 1606
rect 19343 1604 19399 1606
rect 19423 1604 19479 1606
rect 19503 1604 19559 1606
rect 19263 570 19319 572
rect 19343 570 19399 572
rect 19423 570 19479 572
rect 19503 570 19559 572
rect 19263 518 19309 570
rect 19309 518 19319 570
rect 19343 518 19373 570
rect 19373 518 19385 570
rect 19385 518 19399 570
rect 19423 518 19437 570
rect 19437 518 19449 570
rect 19449 518 19479 570
rect 19503 518 19513 570
rect 19513 518 19559 570
rect 19263 516 19319 518
rect 19343 516 19399 518
rect 19423 516 19479 518
rect 19503 516 19559 518
<< metal3 >>
rect 5108 19072 5424 19073
rect 5108 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5424 19072
rect 5108 19007 5424 19008
rect 9823 19072 10139 19073
rect 9823 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10139 19072
rect 9823 19007 10139 19008
rect 14538 19072 14854 19073
rect 14538 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14854 19072
rect 14538 19007 14854 19008
rect 19253 19072 19569 19073
rect 19253 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19569 19072
rect 19253 19007 19569 19008
rect 2751 18528 3067 18529
rect 2751 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3067 18528
rect 2751 18463 3067 18464
rect 7466 18528 7782 18529
rect 7466 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7782 18528
rect 7466 18463 7782 18464
rect 12181 18528 12497 18529
rect 12181 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12497 18528
rect 12181 18463 12497 18464
rect 16896 18528 17212 18529
rect 16896 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17212 18528
rect 16896 18463 17212 18464
rect 5108 17984 5424 17985
rect 5108 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5424 17984
rect 5108 17919 5424 17920
rect 9823 17984 10139 17985
rect 9823 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10139 17984
rect 9823 17919 10139 17920
rect 14538 17984 14854 17985
rect 14538 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14854 17984
rect 14538 17919 14854 17920
rect 19253 17984 19569 17985
rect 19253 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19569 17984
rect 19253 17919 19569 17920
rect 2751 17440 3067 17441
rect 2751 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3067 17440
rect 2751 17375 3067 17376
rect 7466 17440 7782 17441
rect 7466 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7782 17440
rect 7466 17375 7782 17376
rect 12181 17440 12497 17441
rect 12181 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12497 17440
rect 12181 17375 12497 17376
rect 16896 17440 17212 17441
rect 16896 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17212 17440
rect 16896 17375 17212 17376
rect 5108 16896 5424 16897
rect 5108 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5424 16896
rect 5108 16831 5424 16832
rect 9823 16896 10139 16897
rect 9823 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10139 16896
rect 9823 16831 10139 16832
rect 14538 16896 14854 16897
rect 14538 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14854 16896
rect 14538 16831 14854 16832
rect 19253 16896 19569 16897
rect 19253 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19569 16896
rect 19253 16831 19569 16832
rect 6177 16690 6243 16693
rect 8845 16690 8911 16693
rect 6177 16688 8911 16690
rect 6177 16632 6182 16688
rect 6238 16632 8850 16688
rect 8906 16632 8911 16688
rect 6177 16630 8911 16632
rect 6177 16627 6243 16630
rect 8845 16627 8911 16630
rect 9949 16690 10015 16693
rect 10358 16690 10364 16692
rect 9949 16688 10364 16690
rect 9949 16632 9954 16688
rect 10010 16632 10364 16688
rect 9949 16630 10364 16632
rect 9949 16627 10015 16630
rect 10358 16628 10364 16630
rect 10428 16628 10434 16692
rect 2751 16352 3067 16353
rect 2751 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3067 16352
rect 2751 16287 3067 16288
rect 7466 16352 7782 16353
rect 7466 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7782 16352
rect 7466 16287 7782 16288
rect 12181 16352 12497 16353
rect 12181 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12497 16352
rect 12181 16287 12497 16288
rect 16896 16352 17212 16353
rect 16896 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17212 16352
rect 16896 16287 17212 16288
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 19057 16010 19123 16013
rect 17972 16008 19123 16010
rect 17972 15952 19062 16008
rect 19118 15952 19123 16008
rect 17972 15950 19123 15952
rect 17972 15948 17978 15950
rect 19057 15947 19123 15950
rect 5108 15808 5424 15809
rect 5108 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5424 15808
rect 5108 15743 5424 15744
rect 9823 15808 10139 15809
rect 9823 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10139 15808
rect 9823 15743 10139 15744
rect 14538 15808 14854 15809
rect 14538 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14854 15808
rect 14538 15743 14854 15744
rect 19253 15808 19569 15809
rect 19253 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19569 15808
rect 19253 15743 19569 15744
rect 8661 15468 8727 15469
rect 8661 15466 8708 15468
rect 8616 15464 8708 15466
rect 8616 15408 8666 15464
rect 8616 15406 8708 15408
rect 8661 15404 8708 15406
rect 8772 15404 8778 15468
rect 8661 15403 8727 15404
rect 2751 15264 3067 15265
rect 2751 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3067 15264
rect 2751 15199 3067 15200
rect 7466 15264 7782 15265
rect 7466 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7782 15264
rect 7466 15199 7782 15200
rect 12181 15264 12497 15265
rect 12181 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12497 15264
rect 12181 15199 12497 15200
rect 16896 15264 17212 15265
rect 16896 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17212 15264
rect 16896 15199 17212 15200
rect 5108 14720 5424 14721
rect 5108 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5424 14720
rect 5108 14655 5424 14656
rect 9823 14720 10139 14721
rect 9823 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10139 14720
rect 9823 14655 10139 14656
rect 14538 14720 14854 14721
rect 14538 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14854 14720
rect 14538 14655 14854 14656
rect 19253 14720 19569 14721
rect 19253 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19569 14720
rect 19253 14655 19569 14656
rect 2751 14176 3067 14177
rect 2751 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3067 14176
rect 2751 14111 3067 14112
rect 7466 14176 7782 14177
rect 7466 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7782 14176
rect 7466 14111 7782 14112
rect 12181 14176 12497 14177
rect 12181 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12497 14176
rect 12181 14111 12497 14112
rect 16896 14176 17212 14177
rect 16896 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17212 14176
rect 16896 14111 17212 14112
rect 5108 13632 5424 13633
rect 5108 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5424 13632
rect 5108 13567 5424 13568
rect 9823 13632 10139 13633
rect 9823 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10139 13632
rect 9823 13567 10139 13568
rect 14538 13632 14854 13633
rect 14538 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14854 13632
rect 14538 13567 14854 13568
rect 19253 13632 19569 13633
rect 19253 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19569 13632
rect 19253 13567 19569 13568
rect 2751 13088 3067 13089
rect 2751 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3067 13088
rect 2751 13023 3067 13024
rect 7466 13088 7782 13089
rect 7466 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7782 13088
rect 7466 13023 7782 13024
rect 12181 13088 12497 13089
rect 12181 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12497 13088
rect 12181 13023 12497 13024
rect 16896 13088 17212 13089
rect 16896 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17212 13088
rect 16896 13023 17212 13024
rect 6913 12746 6979 12749
rect 8702 12746 8708 12748
rect 6913 12744 8708 12746
rect 6913 12688 6918 12744
rect 6974 12688 8708 12744
rect 6913 12686 8708 12688
rect 6913 12683 6979 12686
rect 8702 12684 8708 12686
rect 8772 12746 8778 12748
rect 9581 12746 9647 12749
rect 11513 12746 11579 12749
rect 8772 12744 11579 12746
rect 8772 12688 9586 12744
rect 9642 12688 11518 12744
rect 11574 12688 11579 12744
rect 8772 12686 11579 12688
rect 8772 12684 8778 12686
rect 9581 12683 9647 12686
rect 11513 12683 11579 12686
rect 5108 12544 5424 12545
rect 5108 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5424 12544
rect 5108 12479 5424 12480
rect 9823 12544 10139 12545
rect 9823 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10139 12544
rect 9823 12479 10139 12480
rect 14538 12544 14854 12545
rect 14538 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14854 12544
rect 14538 12479 14854 12480
rect 19253 12544 19569 12545
rect 19253 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19569 12544
rect 19253 12479 19569 12480
rect 2751 12000 3067 12001
rect 2751 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3067 12000
rect 2751 11935 3067 11936
rect 7466 12000 7782 12001
rect 7466 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7782 12000
rect 7466 11935 7782 11936
rect 12181 12000 12497 12001
rect 12181 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12497 12000
rect 12181 11935 12497 11936
rect 16896 12000 17212 12001
rect 16896 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17212 12000
rect 16896 11935 17212 11936
rect 10593 11794 10659 11797
rect 17902 11794 17908 11796
rect 10593 11792 17908 11794
rect 10593 11736 10598 11792
rect 10654 11736 17908 11792
rect 10593 11734 17908 11736
rect 10593 11731 10659 11734
rect 17902 11732 17908 11734
rect 17972 11732 17978 11796
rect 5108 11456 5424 11457
rect 5108 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5424 11456
rect 5108 11391 5424 11392
rect 9823 11456 10139 11457
rect 9823 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10139 11456
rect 9823 11391 10139 11392
rect 14538 11456 14854 11457
rect 14538 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14854 11456
rect 14538 11391 14854 11392
rect 19253 11456 19569 11457
rect 19253 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19569 11456
rect 19253 11391 19569 11392
rect 2751 10912 3067 10913
rect 2751 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3067 10912
rect 2751 10847 3067 10848
rect 7466 10912 7782 10913
rect 7466 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7782 10912
rect 7466 10847 7782 10848
rect 12181 10912 12497 10913
rect 12181 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12497 10912
rect 12181 10847 12497 10848
rect 16896 10912 17212 10913
rect 16896 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17212 10912
rect 16896 10847 17212 10848
rect 5108 10368 5424 10369
rect 5108 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5424 10368
rect 5108 10303 5424 10304
rect 9823 10368 10139 10369
rect 9823 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10139 10368
rect 9823 10303 10139 10304
rect 14538 10368 14854 10369
rect 14538 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14854 10368
rect 14538 10303 14854 10304
rect 19253 10368 19569 10369
rect 19253 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19569 10368
rect 19253 10303 19569 10304
rect 13629 10298 13695 10301
rect 14365 10298 14431 10301
rect 13629 10296 14431 10298
rect 13629 10240 13634 10296
rect 13690 10240 14370 10296
rect 14426 10240 14431 10296
rect 13629 10238 14431 10240
rect 13629 10235 13695 10238
rect 14365 10235 14431 10238
rect 13077 10162 13143 10165
rect 14181 10162 14247 10165
rect 13077 10160 14247 10162
rect 13077 10104 13082 10160
rect 13138 10104 14186 10160
rect 14242 10104 14247 10160
rect 13077 10102 14247 10104
rect 13077 10099 13143 10102
rect 14181 10099 14247 10102
rect 13629 10026 13695 10029
rect 14733 10026 14799 10029
rect 13629 10024 14799 10026
rect 13629 9968 13634 10024
rect 13690 9968 14738 10024
rect 14794 9968 14799 10024
rect 13629 9966 14799 9968
rect 13629 9963 13695 9966
rect 14733 9963 14799 9966
rect 2751 9824 3067 9825
rect 2751 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3067 9824
rect 2751 9759 3067 9760
rect 7466 9824 7782 9825
rect 7466 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7782 9824
rect 7466 9759 7782 9760
rect 12181 9824 12497 9825
rect 12181 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12497 9824
rect 12181 9759 12497 9760
rect 16896 9824 17212 9825
rect 16896 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17212 9824
rect 16896 9759 17212 9760
rect 10041 9618 10107 9621
rect 10777 9618 10843 9621
rect 10041 9616 10843 9618
rect 10041 9560 10046 9616
rect 10102 9560 10782 9616
rect 10838 9560 10843 9616
rect 10041 9558 10843 9560
rect 10041 9555 10107 9558
rect 10777 9555 10843 9558
rect 5108 9280 5424 9281
rect 5108 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5424 9280
rect 5108 9215 5424 9216
rect 9823 9280 10139 9281
rect 9823 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10139 9280
rect 9823 9215 10139 9216
rect 14538 9280 14854 9281
rect 14538 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14854 9280
rect 14538 9215 14854 9216
rect 19253 9280 19569 9281
rect 19253 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19569 9280
rect 19253 9215 19569 9216
rect 2751 8736 3067 8737
rect 2751 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3067 8736
rect 2751 8671 3067 8672
rect 7466 8736 7782 8737
rect 7466 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7782 8736
rect 7466 8671 7782 8672
rect 12181 8736 12497 8737
rect 12181 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12497 8736
rect 12181 8671 12497 8672
rect 16896 8736 17212 8737
rect 16896 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17212 8736
rect 16896 8671 17212 8672
rect 5108 8192 5424 8193
rect 5108 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5424 8192
rect 5108 8127 5424 8128
rect 9823 8192 10139 8193
rect 9823 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10139 8192
rect 9823 8127 10139 8128
rect 14538 8192 14854 8193
rect 14538 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14854 8192
rect 14538 8127 14854 8128
rect 19253 8192 19569 8193
rect 19253 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19569 8192
rect 19253 8127 19569 8128
rect 2751 7648 3067 7649
rect 2751 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3067 7648
rect 2751 7583 3067 7584
rect 7466 7648 7782 7649
rect 7466 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7782 7648
rect 7466 7583 7782 7584
rect 12181 7648 12497 7649
rect 12181 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12497 7648
rect 12181 7583 12497 7584
rect 16896 7648 17212 7649
rect 16896 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17212 7648
rect 16896 7583 17212 7584
rect 5108 7104 5424 7105
rect 5108 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5424 7104
rect 5108 7039 5424 7040
rect 9823 7104 10139 7105
rect 9823 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10139 7104
rect 9823 7039 10139 7040
rect 14538 7104 14854 7105
rect 14538 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14854 7104
rect 14538 7039 14854 7040
rect 19253 7104 19569 7105
rect 19253 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19569 7104
rect 19253 7039 19569 7040
rect 10358 6836 10364 6900
rect 10428 6898 10434 6900
rect 11145 6898 11211 6901
rect 10428 6896 11211 6898
rect 10428 6840 11150 6896
rect 11206 6840 11211 6896
rect 10428 6838 11211 6840
rect 10428 6836 10434 6838
rect 11145 6835 11211 6838
rect 2751 6560 3067 6561
rect 2751 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3067 6560
rect 2751 6495 3067 6496
rect 7466 6560 7782 6561
rect 7466 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7782 6560
rect 7466 6495 7782 6496
rect 12181 6560 12497 6561
rect 12181 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12497 6560
rect 12181 6495 12497 6496
rect 16896 6560 17212 6561
rect 16896 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17212 6560
rect 16896 6495 17212 6496
rect 5108 6016 5424 6017
rect 5108 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5424 6016
rect 5108 5951 5424 5952
rect 9823 6016 10139 6017
rect 9823 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10139 6016
rect 9823 5951 10139 5952
rect 14538 6016 14854 6017
rect 14538 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14854 6016
rect 14538 5951 14854 5952
rect 19253 6016 19569 6017
rect 19253 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19569 6016
rect 19253 5951 19569 5952
rect 2751 5472 3067 5473
rect 2751 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3067 5472
rect 2751 5407 3067 5408
rect 7466 5472 7782 5473
rect 7466 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7782 5472
rect 7466 5407 7782 5408
rect 12181 5472 12497 5473
rect 12181 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12497 5472
rect 12181 5407 12497 5408
rect 16896 5472 17212 5473
rect 16896 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17212 5472
rect 16896 5407 17212 5408
rect 5108 4928 5424 4929
rect 5108 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5424 4928
rect 5108 4863 5424 4864
rect 9823 4928 10139 4929
rect 9823 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10139 4928
rect 9823 4863 10139 4864
rect 14538 4928 14854 4929
rect 14538 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14854 4928
rect 14538 4863 14854 4864
rect 19253 4928 19569 4929
rect 19253 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19569 4928
rect 19253 4863 19569 4864
rect 2751 4384 3067 4385
rect 2751 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3067 4384
rect 2751 4319 3067 4320
rect 7466 4384 7782 4385
rect 7466 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7782 4384
rect 7466 4319 7782 4320
rect 12181 4384 12497 4385
rect 12181 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12497 4384
rect 12181 4319 12497 4320
rect 16896 4384 17212 4385
rect 16896 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17212 4384
rect 16896 4319 17212 4320
rect 5108 3840 5424 3841
rect 5108 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5424 3840
rect 5108 3775 5424 3776
rect 9823 3840 10139 3841
rect 9823 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10139 3840
rect 9823 3775 10139 3776
rect 14538 3840 14854 3841
rect 14538 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14854 3840
rect 14538 3775 14854 3776
rect 19253 3840 19569 3841
rect 19253 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19569 3840
rect 19253 3775 19569 3776
rect 2751 3296 3067 3297
rect 2751 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3067 3296
rect 2751 3231 3067 3232
rect 7466 3296 7782 3297
rect 7466 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7782 3296
rect 7466 3231 7782 3232
rect 12181 3296 12497 3297
rect 12181 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12497 3296
rect 12181 3231 12497 3232
rect 16896 3296 17212 3297
rect 16896 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17212 3296
rect 16896 3231 17212 3232
rect 5108 2752 5424 2753
rect 5108 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5424 2752
rect 5108 2687 5424 2688
rect 9823 2752 10139 2753
rect 9823 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10139 2752
rect 9823 2687 10139 2688
rect 14538 2752 14854 2753
rect 14538 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14854 2752
rect 14538 2687 14854 2688
rect 19253 2752 19569 2753
rect 19253 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19569 2752
rect 19253 2687 19569 2688
rect 2751 2208 3067 2209
rect 2751 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3067 2208
rect 2751 2143 3067 2144
rect 7466 2208 7782 2209
rect 7466 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7782 2208
rect 7466 2143 7782 2144
rect 12181 2208 12497 2209
rect 12181 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12497 2208
rect 12181 2143 12497 2144
rect 16896 2208 17212 2209
rect 16896 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17212 2208
rect 16896 2143 17212 2144
rect 5108 1664 5424 1665
rect 5108 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5424 1664
rect 5108 1599 5424 1600
rect 9823 1664 10139 1665
rect 9823 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10139 1664
rect 9823 1599 10139 1600
rect 14538 1664 14854 1665
rect 14538 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14854 1664
rect 14538 1599 14854 1600
rect 19253 1664 19569 1665
rect 19253 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19569 1664
rect 19253 1599 19569 1600
rect 2751 1120 3067 1121
rect 2751 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3067 1120
rect 2751 1055 3067 1056
rect 7466 1120 7782 1121
rect 7466 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7782 1120
rect 7466 1055 7782 1056
rect 12181 1120 12497 1121
rect 12181 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12497 1120
rect 12181 1055 12497 1056
rect 16896 1120 17212 1121
rect 16896 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17212 1120
rect 16896 1055 17212 1056
rect 5108 576 5424 577
rect 5108 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5424 576
rect 5108 511 5424 512
rect 9823 576 10139 577
rect 9823 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10139 576
rect 9823 511 10139 512
rect 14538 576 14854 577
rect 14538 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14854 576
rect 14538 511 14854 512
rect 19253 576 19569 577
rect 19253 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19569 576
rect 19253 511 19569 512
<< via3 >>
rect 5114 19068 5178 19072
rect 5114 19012 5118 19068
rect 5118 19012 5174 19068
rect 5174 19012 5178 19068
rect 5114 19008 5178 19012
rect 5194 19068 5258 19072
rect 5194 19012 5198 19068
rect 5198 19012 5254 19068
rect 5254 19012 5258 19068
rect 5194 19008 5258 19012
rect 5274 19068 5338 19072
rect 5274 19012 5278 19068
rect 5278 19012 5334 19068
rect 5334 19012 5338 19068
rect 5274 19008 5338 19012
rect 5354 19068 5418 19072
rect 5354 19012 5358 19068
rect 5358 19012 5414 19068
rect 5414 19012 5418 19068
rect 5354 19008 5418 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 10069 19068 10133 19072
rect 10069 19012 10073 19068
rect 10073 19012 10129 19068
rect 10129 19012 10133 19068
rect 10069 19008 10133 19012
rect 14544 19068 14608 19072
rect 14544 19012 14548 19068
rect 14548 19012 14604 19068
rect 14604 19012 14608 19068
rect 14544 19008 14608 19012
rect 14624 19068 14688 19072
rect 14624 19012 14628 19068
rect 14628 19012 14684 19068
rect 14684 19012 14688 19068
rect 14624 19008 14688 19012
rect 14704 19068 14768 19072
rect 14704 19012 14708 19068
rect 14708 19012 14764 19068
rect 14764 19012 14768 19068
rect 14704 19008 14768 19012
rect 14784 19068 14848 19072
rect 14784 19012 14788 19068
rect 14788 19012 14844 19068
rect 14844 19012 14848 19068
rect 14784 19008 14848 19012
rect 19259 19068 19323 19072
rect 19259 19012 19263 19068
rect 19263 19012 19319 19068
rect 19319 19012 19323 19068
rect 19259 19008 19323 19012
rect 19339 19068 19403 19072
rect 19339 19012 19343 19068
rect 19343 19012 19399 19068
rect 19399 19012 19403 19068
rect 19339 19008 19403 19012
rect 19419 19068 19483 19072
rect 19419 19012 19423 19068
rect 19423 19012 19479 19068
rect 19479 19012 19483 19068
rect 19419 19008 19483 19012
rect 19499 19068 19563 19072
rect 19499 19012 19503 19068
rect 19503 19012 19559 19068
rect 19559 19012 19563 19068
rect 19499 19008 19563 19012
rect 2757 18524 2821 18528
rect 2757 18468 2761 18524
rect 2761 18468 2817 18524
rect 2817 18468 2821 18524
rect 2757 18464 2821 18468
rect 2837 18524 2901 18528
rect 2837 18468 2841 18524
rect 2841 18468 2897 18524
rect 2897 18468 2901 18524
rect 2837 18464 2901 18468
rect 2917 18524 2981 18528
rect 2917 18468 2921 18524
rect 2921 18468 2977 18524
rect 2977 18468 2981 18524
rect 2917 18464 2981 18468
rect 2997 18524 3061 18528
rect 2997 18468 3001 18524
rect 3001 18468 3057 18524
rect 3057 18468 3061 18524
rect 2997 18464 3061 18468
rect 7472 18524 7536 18528
rect 7472 18468 7476 18524
rect 7476 18468 7532 18524
rect 7532 18468 7536 18524
rect 7472 18464 7536 18468
rect 7552 18524 7616 18528
rect 7552 18468 7556 18524
rect 7556 18468 7612 18524
rect 7612 18468 7616 18524
rect 7552 18464 7616 18468
rect 7632 18524 7696 18528
rect 7632 18468 7636 18524
rect 7636 18468 7692 18524
rect 7692 18468 7696 18524
rect 7632 18464 7696 18468
rect 7712 18524 7776 18528
rect 7712 18468 7716 18524
rect 7716 18468 7772 18524
rect 7772 18468 7776 18524
rect 7712 18464 7776 18468
rect 12187 18524 12251 18528
rect 12187 18468 12191 18524
rect 12191 18468 12247 18524
rect 12247 18468 12251 18524
rect 12187 18464 12251 18468
rect 12267 18524 12331 18528
rect 12267 18468 12271 18524
rect 12271 18468 12327 18524
rect 12327 18468 12331 18524
rect 12267 18464 12331 18468
rect 12347 18524 12411 18528
rect 12347 18468 12351 18524
rect 12351 18468 12407 18524
rect 12407 18468 12411 18524
rect 12347 18464 12411 18468
rect 12427 18524 12491 18528
rect 12427 18468 12431 18524
rect 12431 18468 12487 18524
rect 12487 18468 12491 18524
rect 12427 18464 12491 18468
rect 16902 18524 16966 18528
rect 16902 18468 16906 18524
rect 16906 18468 16962 18524
rect 16962 18468 16966 18524
rect 16902 18464 16966 18468
rect 16982 18524 17046 18528
rect 16982 18468 16986 18524
rect 16986 18468 17042 18524
rect 17042 18468 17046 18524
rect 16982 18464 17046 18468
rect 17062 18524 17126 18528
rect 17062 18468 17066 18524
rect 17066 18468 17122 18524
rect 17122 18468 17126 18524
rect 17062 18464 17126 18468
rect 17142 18524 17206 18528
rect 17142 18468 17146 18524
rect 17146 18468 17202 18524
rect 17202 18468 17206 18524
rect 17142 18464 17206 18468
rect 5114 17980 5178 17984
rect 5114 17924 5118 17980
rect 5118 17924 5174 17980
rect 5174 17924 5178 17980
rect 5114 17920 5178 17924
rect 5194 17980 5258 17984
rect 5194 17924 5198 17980
rect 5198 17924 5254 17980
rect 5254 17924 5258 17980
rect 5194 17920 5258 17924
rect 5274 17980 5338 17984
rect 5274 17924 5278 17980
rect 5278 17924 5334 17980
rect 5334 17924 5338 17980
rect 5274 17920 5338 17924
rect 5354 17980 5418 17984
rect 5354 17924 5358 17980
rect 5358 17924 5414 17980
rect 5414 17924 5418 17980
rect 5354 17920 5418 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 10069 17980 10133 17984
rect 10069 17924 10073 17980
rect 10073 17924 10129 17980
rect 10129 17924 10133 17980
rect 10069 17920 10133 17924
rect 14544 17980 14608 17984
rect 14544 17924 14548 17980
rect 14548 17924 14604 17980
rect 14604 17924 14608 17980
rect 14544 17920 14608 17924
rect 14624 17980 14688 17984
rect 14624 17924 14628 17980
rect 14628 17924 14684 17980
rect 14684 17924 14688 17980
rect 14624 17920 14688 17924
rect 14704 17980 14768 17984
rect 14704 17924 14708 17980
rect 14708 17924 14764 17980
rect 14764 17924 14768 17980
rect 14704 17920 14768 17924
rect 14784 17980 14848 17984
rect 14784 17924 14788 17980
rect 14788 17924 14844 17980
rect 14844 17924 14848 17980
rect 14784 17920 14848 17924
rect 19259 17980 19323 17984
rect 19259 17924 19263 17980
rect 19263 17924 19319 17980
rect 19319 17924 19323 17980
rect 19259 17920 19323 17924
rect 19339 17980 19403 17984
rect 19339 17924 19343 17980
rect 19343 17924 19399 17980
rect 19399 17924 19403 17980
rect 19339 17920 19403 17924
rect 19419 17980 19483 17984
rect 19419 17924 19423 17980
rect 19423 17924 19479 17980
rect 19479 17924 19483 17980
rect 19419 17920 19483 17924
rect 19499 17980 19563 17984
rect 19499 17924 19503 17980
rect 19503 17924 19559 17980
rect 19559 17924 19563 17980
rect 19499 17920 19563 17924
rect 2757 17436 2821 17440
rect 2757 17380 2761 17436
rect 2761 17380 2817 17436
rect 2817 17380 2821 17436
rect 2757 17376 2821 17380
rect 2837 17436 2901 17440
rect 2837 17380 2841 17436
rect 2841 17380 2897 17436
rect 2897 17380 2901 17436
rect 2837 17376 2901 17380
rect 2917 17436 2981 17440
rect 2917 17380 2921 17436
rect 2921 17380 2977 17436
rect 2977 17380 2981 17436
rect 2917 17376 2981 17380
rect 2997 17436 3061 17440
rect 2997 17380 3001 17436
rect 3001 17380 3057 17436
rect 3057 17380 3061 17436
rect 2997 17376 3061 17380
rect 7472 17436 7536 17440
rect 7472 17380 7476 17436
rect 7476 17380 7532 17436
rect 7532 17380 7536 17436
rect 7472 17376 7536 17380
rect 7552 17436 7616 17440
rect 7552 17380 7556 17436
rect 7556 17380 7612 17436
rect 7612 17380 7616 17436
rect 7552 17376 7616 17380
rect 7632 17436 7696 17440
rect 7632 17380 7636 17436
rect 7636 17380 7692 17436
rect 7692 17380 7696 17436
rect 7632 17376 7696 17380
rect 7712 17436 7776 17440
rect 7712 17380 7716 17436
rect 7716 17380 7772 17436
rect 7772 17380 7776 17436
rect 7712 17376 7776 17380
rect 12187 17436 12251 17440
rect 12187 17380 12191 17436
rect 12191 17380 12247 17436
rect 12247 17380 12251 17436
rect 12187 17376 12251 17380
rect 12267 17436 12331 17440
rect 12267 17380 12271 17436
rect 12271 17380 12327 17436
rect 12327 17380 12331 17436
rect 12267 17376 12331 17380
rect 12347 17436 12411 17440
rect 12347 17380 12351 17436
rect 12351 17380 12407 17436
rect 12407 17380 12411 17436
rect 12347 17376 12411 17380
rect 12427 17436 12491 17440
rect 12427 17380 12431 17436
rect 12431 17380 12487 17436
rect 12487 17380 12491 17436
rect 12427 17376 12491 17380
rect 16902 17436 16966 17440
rect 16902 17380 16906 17436
rect 16906 17380 16962 17436
rect 16962 17380 16966 17436
rect 16902 17376 16966 17380
rect 16982 17436 17046 17440
rect 16982 17380 16986 17436
rect 16986 17380 17042 17436
rect 17042 17380 17046 17436
rect 16982 17376 17046 17380
rect 17062 17436 17126 17440
rect 17062 17380 17066 17436
rect 17066 17380 17122 17436
rect 17122 17380 17126 17436
rect 17062 17376 17126 17380
rect 17142 17436 17206 17440
rect 17142 17380 17146 17436
rect 17146 17380 17202 17436
rect 17202 17380 17206 17436
rect 17142 17376 17206 17380
rect 5114 16892 5178 16896
rect 5114 16836 5118 16892
rect 5118 16836 5174 16892
rect 5174 16836 5178 16892
rect 5114 16832 5178 16836
rect 5194 16892 5258 16896
rect 5194 16836 5198 16892
rect 5198 16836 5254 16892
rect 5254 16836 5258 16892
rect 5194 16832 5258 16836
rect 5274 16892 5338 16896
rect 5274 16836 5278 16892
rect 5278 16836 5334 16892
rect 5334 16836 5338 16892
rect 5274 16832 5338 16836
rect 5354 16892 5418 16896
rect 5354 16836 5358 16892
rect 5358 16836 5414 16892
rect 5414 16836 5418 16892
rect 5354 16832 5418 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 10069 16892 10133 16896
rect 10069 16836 10073 16892
rect 10073 16836 10129 16892
rect 10129 16836 10133 16892
rect 10069 16832 10133 16836
rect 14544 16892 14608 16896
rect 14544 16836 14548 16892
rect 14548 16836 14604 16892
rect 14604 16836 14608 16892
rect 14544 16832 14608 16836
rect 14624 16892 14688 16896
rect 14624 16836 14628 16892
rect 14628 16836 14684 16892
rect 14684 16836 14688 16892
rect 14624 16832 14688 16836
rect 14704 16892 14768 16896
rect 14704 16836 14708 16892
rect 14708 16836 14764 16892
rect 14764 16836 14768 16892
rect 14704 16832 14768 16836
rect 14784 16892 14848 16896
rect 14784 16836 14788 16892
rect 14788 16836 14844 16892
rect 14844 16836 14848 16892
rect 14784 16832 14848 16836
rect 19259 16892 19323 16896
rect 19259 16836 19263 16892
rect 19263 16836 19319 16892
rect 19319 16836 19323 16892
rect 19259 16832 19323 16836
rect 19339 16892 19403 16896
rect 19339 16836 19343 16892
rect 19343 16836 19399 16892
rect 19399 16836 19403 16892
rect 19339 16832 19403 16836
rect 19419 16892 19483 16896
rect 19419 16836 19423 16892
rect 19423 16836 19479 16892
rect 19479 16836 19483 16892
rect 19419 16832 19483 16836
rect 19499 16892 19563 16896
rect 19499 16836 19503 16892
rect 19503 16836 19559 16892
rect 19559 16836 19563 16892
rect 19499 16832 19563 16836
rect 10364 16628 10428 16692
rect 2757 16348 2821 16352
rect 2757 16292 2761 16348
rect 2761 16292 2817 16348
rect 2817 16292 2821 16348
rect 2757 16288 2821 16292
rect 2837 16348 2901 16352
rect 2837 16292 2841 16348
rect 2841 16292 2897 16348
rect 2897 16292 2901 16348
rect 2837 16288 2901 16292
rect 2917 16348 2981 16352
rect 2917 16292 2921 16348
rect 2921 16292 2977 16348
rect 2977 16292 2981 16348
rect 2917 16288 2981 16292
rect 2997 16348 3061 16352
rect 2997 16292 3001 16348
rect 3001 16292 3057 16348
rect 3057 16292 3061 16348
rect 2997 16288 3061 16292
rect 7472 16348 7536 16352
rect 7472 16292 7476 16348
rect 7476 16292 7532 16348
rect 7532 16292 7536 16348
rect 7472 16288 7536 16292
rect 7552 16348 7616 16352
rect 7552 16292 7556 16348
rect 7556 16292 7612 16348
rect 7612 16292 7616 16348
rect 7552 16288 7616 16292
rect 7632 16348 7696 16352
rect 7632 16292 7636 16348
rect 7636 16292 7692 16348
rect 7692 16292 7696 16348
rect 7632 16288 7696 16292
rect 7712 16348 7776 16352
rect 7712 16292 7716 16348
rect 7716 16292 7772 16348
rect 7772 16292 7776 16348
rect 7712 16288 7776 16292
rect 12187 16348 12251 16352
rect 12187 16292 12191 16348
rect 12191 16292 12247 16348
rect 12247 16292 12251 16348
rect 12187 16288 12251 16292
rect 12267 16348 12331 16352
rect 12267 16292 12271 16348
rect 12271 16292 12327 16348
rect 12327 16292 12331 16348
rect 12267 16288 12331 16292
rect 12347 16348 12411 16352
rect 12347 16292 12351 16348
rect 12351 16292 12407 16348
rect 12407 16292 12411 16348
rect 12347 16288 12411 16292
rect 12427 16348 12491 16352
rect 12427 16292 12431 16348
rect 12431 16292 12487 16348
rect 12487 16292 12491 16348
rect 12427 16288 12491 16292
rect 16902 16348 16966 16352
rect 16902 16292 16906 16348
rect 16906 16292 16962 16348
rect 16962 16292 16966 16348
rect 16902 16288 16966 16292
rect 16982 16348 17046 16352
rect 16982 16292 16986 16348
rect 16986 16292 17042 16348
rect 17042 16292 17046 16348
rect 16982 16288 17046 16292
rect 17062 16348 17126 16352
rect 17062 16292 17066 16348
rect 17066 16292 17122 16348
rect 17122 16292 17126 16348
rect 17062 16288 17126 16292
rect 17142 16348 17206 16352
rect 17142 16292 17146 16348
rect 17146 16292 17202 16348
rect 17202 16292 17206 16348
rect 17142 16288 17206 16292
rect 17908 15948 17972 16012
rect 5114 15804 5178 15808
rect 5114 15748 5118 15804
rect 5118 15748 5174 15804
rect 5174 15748 5178 15804
rect 5114 15744 5178 15748
rect 5194 15804 5258 15808
rect 5194 15748 5198 15804
rect 5198 15748 5254 15804
rect 5254 15748 5258 15804
rect 5194 15744 5258 15748
rect 5274 15804 5338 15808
rect 5274 15748 5278 15804
rect 5278 15748 5334 15804
rect 5334 15748 5338 15804
rect 5274 15744 5338 15748
rect 5354 15804 5418 15808
rect 5354 15748 5358 15804
rect 5358 15748 5414 15804
rect 5414 15748 5418 15804
rect 5354 15744 5418 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 10069 15804 10133 15808
rect 10069 15748 10073 15804
rect 10073 15748 10129 15804
rect 10129 15748 10133 15804
rect 10069 15744 10133 15748
rect 14544 15804 14608 15808
rect 14544 15748 14548 15804
rect 14548 15748 14604 15804
rect 14604 15748 14608 15804
rect 14544 15744 14608 15748
rect 14624 15804 14688 15808
rect 14624 15748 14628 15804
rect 14628 15748 14684 15804
rect 14684 15748 14688 15804
rect 14624 15744 14688 15748
rect 14704 15804 14768 15808
rect 14704 15748 14708 15804
rect 14708 15748 14764 15804
rect 14764 15748 14768 15804
rect 14704 15744 14768 15748
rect 14784 15804 14848 15808
rect 14784 15748 14788 15804
rect 14788 15748 14844 15804
rect 14844 15748 14848 15804
rect 14784 15744 14848 15748
rect 19259 15804 19323 15808
rect 19259 15748 19263 15804
rect 19263 15748 19319 15804
rect 19319 15748 19323 15804
rect 19259 15744 19323 15748
rect 19339 15804 19403 15808
rect 19339 15748 19343 15804
rect 19343 15748 19399 15804
rect 19399 15748 19403 15804
rect 19339 15744 19403 15748
rect 19419 15804 19483 15808
rect 19419 15748 19423 15804
rect 19423 15748 19479 15804
rect 19479 15748 19483 15804
rect 19419 15744 19483 15748
rect 19499 15804 19563 15808
rect 19499 15748 19503 15804
rect 19503 15748 19559 15804
rect 19559 15748 19563 15804
rect 19499 15744 19563 15748
rect 8708 15464 8772 15468
rect 8708 15408 8722 15464
rect 8722 15408 8772 15464
rect 8708 15404 8772 15408
rect 2757 15260 2821 15264
rect 2757 15204 2761 15260
rect 2761 15204 2817 15260
rect 2817 15204 2821 15260
rect 2757 15200 2821 15204
rect 2837 15260 2901 15264
rect 2837 15204 2841 15260
rect 2841 15204 2897 15260
rect 2897 15204 2901 15260
rect 2837 15200 2901 15204
rect 2917 15260 2981 15264
rect 2917 15204 2921 15260
rect 2921 15204 2977 15260
rect 2977 15204 2981 15260
rect 2917 15200 2981 15204
rect 2997 15260 3061 15264
rect 2997 15204 3001 15260
rect 3001 15204 3057 15260
rect 3057 15204 3061 15260
rect 2997 15200 3061 15204
rect 7472 15260 7536 15264
rect 7472 15204 7476 15260
rect 7476 15204 7532 15260
rect 7532 15204 7536 15260
rect 7472 15200 7536 15204
rect 7552 15260 7616 15264
rect 7552 15204 7556 15260
rect 7556 15204 7612 15260
rect 7612 15204 7616 15260
rect 7552 15200 7616 15204
rect 7632 15260 7696 15264
rect 7632 15204 7636 15260
rect 7636 15204 7692 15260
rect 7692 15204 7696 15260
rect 7632 15200 7696 15204
rect 7712 15260 7776 15264
rect 7712 15204 7716 15260
rect 7716 15204 7772 15260
rect 7772 15204 7776 15260
rect 7712 15200 7776 15204
rect 12187 15260 12251 15264
rect 12187 15204 12191 15260
rect 12191 15204 12247 15260
rect 12247 15204 12251 15260
rect 12187 15200 12251 15204
rect 12267 15260 12331 15264
rect 12267 15204 12271 15260
rect 12271 15204 12327 15260
rect 12327 15204 12331 15260
rect 12267 15200 12331 15204
rect 12347 15260 12411 15264
rect 12347 15204 12351 15260
rect 12351 15204 12407 15260
rect 12407 15204 12411 15260
rect 12347 15200 12411 15204
rect 12427 15260 12491 15264
rect 12427 15204 12431 15260
rect 12431 15204 12487 15260
rect 12487 15204 12491 15260
rect 12427 15200 12491 15204
rect 16902 15260 16966 15264
rect 16902 15204 16906 15260
rect 16906 15204 16962 15260
rect 16962 15204 16966 15260
rect 16902 15200 16966 15204
rect 16982 15260 17046 15264
rect 16982 15204 16986 15260
rect 16986 15204 17042 15260
rect 17042 15204 17046 15260
rect 16982 15200 17046 15204
rect 17062 15260 17126 15264
rect 17062 15204 17066 15260
rect 17066 15204 17122 15260
rect 17122 15204 17126 15260
rect 17062 15200 17126 15204
rect 17142 15260 17206 15264
rect 17142 15204 17146 15260
rect 17146 15204 17202 15260
rect 17202 15204 17206 15260
rect 17142 15200 17206 15204
rect 5114 14716 5178 14720
rect 5114 14660 5118 14716
rect 5118 14660 5174 14716
rect 5174 14660 5178 14716
rect 5114 14656 5178 14660
rect 5194 14716 5258 14720
rect 5194 14660 5198 14716
rect 5198 14660 5254 14716
rect 5254 14660 5258 14716
rect 5194 14656 5258 14660
rect 5274 14716 5338 14720
rect 5274 14660 5278 14716
rect 5278 14660 5334 14716
rect 5334 14660 5338 14716
rect 5274 14656 5338 14660
rect 5354 14716 5418 14720
rect 5354 14660 5358 14716
rect 5358 14660 5414 14716
rect 5414 14660 5418 14716
rect 5354 14656 5418 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 10069 14716 10133 14720
rect 10069 14660 10073 14716
rect 10073 14660 10129 14716
rect 10129 14660 10133 14716
rect 10069 14656 10133 14660
rect 14544 14716 14608 14720
rect 14544 14660 14548 14716
rect 14548 14660 14604 14716
rect 14604 14660 14608 14716
rect 14544 14656 14608 14660
rect 14624 14716 14688 14720
rect 14624 14660 14628 14716
rect 14628 14660 14684 14716
rect 14684 14660 14688 14716
rect 14624 14656 14688 14660
rect 14704 14716 14768 14720
rect 14704 14660 14708 14716
rect 14708 14660 14764 14716
rect 14764 14660 14768 14716
rect 14704 14656 14768 14660
rect 14784 14716 14848 14720
rect 14784 14660 14788 14716
rect 14788 14660 14844 14716
rect 14844 14660 14848 14716
rect 14784 14656 14848 14660
rect 19259 14716 19323 14720
rect 19259 14660 19263 14716
rect 19263 14660 19319 14716
rect 19319 14660 19323 14716
rect 19259 14656 19323 14660
rect 19339 14716 19403 14720
rect 19339 14660 19343 14716
rect 19343 14660 19399 14716
rect 19399 14660 19403 14716
rect 19339 14656 19403 14660
rect 19419 14716 19483 14720
rect 19419 14660 19423 14716
rect 19423 14660 19479 14716
rect 19479 14660 19483 14716
rect 19419 14656 19483 14660
rect 19499 14716 19563 14720
rect 19499 14660 19503 14716
rect 19503 14660 19559 14716
rect 19559 14660 19563 14716
rect 19499 14656 19563 14660
rect 2757 14172 2821 14176
rect 2757 14116 2761 14172
rect 2761 14116 2817 14172
rect 2817 14116 2821 14172
rect 2757 14112 2821 14116
rect 2837 14172 2901 14176
rect 2837 14116 2841 14172
rect 2841 14116 2897 14172
rect 2897 14116 2901 14172
rect 2837 14112 2901 14116
rect 2917 14172 2981 14176
rect 2917 14116 2921 14172
rect 2921 14116 2977 14172
rect 2977 14116 2981 14172
rect 2917 14112 2981 14116
rect 2997 14172 3061 14176
rect 2997 14116 3001 14172
rect 3001 14116 3057 14172
rect 3057 14116 3061 14172
rect 2997 14112 3061 14116
rect 7472 14172 7536 14176
rect 7472 14116 7476 14172
rect 7476 14116 7532 14172
rect 7532 14116 7536 14172
rect 7472 14112 7536 14116
rect 7552 14172 7616 14176
rect 7552 14116 7556 14172
rect 7556 14116 7612 14172
rect 7612 14116 7616 14172
rect 7552 14112 7616 14116
rect 7632 14172 7696 14176
rect 7632 14116 7636 14172
rect 7636 14116 7692 14172
rect 7692 14116 7696 14172
rect 7632 14112 7696 14116
rect 7712 14172 7776 14176
rect 7712 14116 7716 14172
rect 7716 14116 7772 14172
rect 7772 14116 7776 14172
rect 7712 14112 7776 14116
rect 12187 14172 12251 14176
rect 12187 14116 12191 14172
rect 12191 14116 12247 14172
rect 12247 14116 12251 14172
rect 12187 14112 12251 14116
rect 12267 14172 12331 14176
rect 12267 14116 12271 14172
rect 12271 14116 12327 14172
rect 12327 14116 12331 14172
rect 12267 14112 12331 14116
rect 12347 14172 12411 14176
rect 12347 14116 12351 14172
rect 12351 14116 12407 14172
rect 12407 14116 12411 14172
rect 12347 14112 12411 14116
rect 12427 14172 12491 14176
rect 12427 14116 12431 14172
rect 12431 14116 12487 14172
rect 12487 14116 12491 14172
rect 12427 14112 12491 14116
rect 16902 14172 16966 14176
rect 16902 14116 16906 14172
rect 16906 14116 16962 14172
rect 16962 14116 16966 14172
rect 16902 14112 16966 14116
rect 16982 14172 17046 14176
rect 16982 14116 16986 14172
rect 16986 14116 17042 14172
rect 17042 14116 17046 14172
rect 16982 14112 17046 14116
rect 17062 14172 17126 14176
rect 17062 14116 17066 14172
rect 17066 14116 17122 14172
rect 17122 14116 17126 14172
rect 17062 14112 17126 14116
rect 17142 14172 17206 14176
rect 17142 14116 17146 14172
rect 17146 14116 17202 14172
rect 17202 14116 17206 14172
rect 17142 14112 17206 14116
rect 5114 13628 5178 13632
rect 5114 13572 5118 13628
rect 5118 13572 5174 13628
rect 5174 13572 5178 13628
rect 5114 13568 5178 13572
rect 5194 13628 5258 13632
rect 5194 13572 5198 13628
rect 5198 13572 5254 13628
rect 5254 13572 5258 13628
rect 5194 13568 5258 13572
rect 5274 13628 5338 13632
rect 5274 13572 5278 13628
rect 5278 13572 5334 13628
rect 5334 13572 5338 13628
rect 5274 13568 5338 13572
rect 5354 13628 5418 13632
rect 5354 13572 5358 13628
rect 5358 13572 5414 13628
rect 5414 13572 5418 13628
rect 5354 13568 5418 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 10069 13628 10133 13632
rect 10069 13572 10073 13628
rect 10073 13572 10129 13628
rect 10129 13572 10133 13628
rect 10069 13568 10133 13572
rect 14544 13628 14608 13632
rect 14544 13572 14548 13628
rect 14548 13572 14604 13628
rect 14604 13572 14608 13628
rect 14544 13568 14608 13572
rect 14624 13628 14688 13632
rect 14624 13572 14628 13628
rect 14628 13572 14684 13628
rect 14684 13572 14688 13628
rect 14624 13568 14688 13572
rect 14704 13628 14768 13632
rect 14704 13572 14708 13628
rect 14708 13572 14764 13628
rect 14764 13572 14768 13628
rect 14704 13568 14768 13572
rect 14784 13628 14848 13632
rect 14784 13572 14788 13628
rect 14788 13572 14844 13628
rect 14844 13572 14848 13628
rect 14784 13568 14848 13572
rect 19259 13628 19323 13632
rect 19259 13572 19263 13628
rect 19263 13572 19319 13628
rect 19319 13572 19323 13628
rect 19259 13568 19323 13572
rect 19339 13628 19403 13632
rect 19339 13572 19343 13628
rect 19343 13572 19399 13628
rect 19399 13572 19403 13628
rect 19339 13568 19403 13572
rect 19419 13628 19483 13632
rect 19419 13572 19423 13628
rect 19423 13572 19479 13628
rect 19479 13572 19483 13628
rect 19419 13568 19483 13572
rect 19499 13628 19563 13632
rect 19499 13572 19503 13628
rect 19503 13572 19559 13628
rect 19559 13572 19563 13628
rect 19499 13568 19563 13572
rect 2757 13084 2821 13088
rect 2757 13028 2761 13084
rect 2761 13028 2817 13084
rect 2817 13028 2821 13084
rect 2757 13024 2821 13028
rect 2837 13084 2901 13088
rect 2837 13028 2841 13084
rect 2841 13028 2897 13084
rect 2897 13028 2901 13084
rect 2837 13024 2901 13028
rect 2917 13084 2981 13088
rect 2917 13028 2921 13084
rect 2921 13028 2977 13084
rect 2977 13028 2981 13084
rect 2917 13024 2981 13028
rect 2997 13084 3061 13088
rect 2997 13028 3001 13084
rect 3001 13028 3057 13084
rect 3057 13028 3061 13084
rect 2997 13024 3061 13028
rect 7472 13084 7536 13088
rect 7472 13028 7476 13084
rect 7476 13028 7532 13084
rect 7532 13028 7536 13084
rect 7472 13024 7536 13028
rect 7552 13084 7616 13088
rect 7552 13028 7556 13084
rect 7556 13028 7612 13084
rect 7612 13028 7616 13084
rect 7552 13024 7616 13028
rect 7632 13084 7696 13088
rect 7632 13028 7636 13084
rect 7636 13028 7692 13084
rect 7692 13028 7696 13084
rect 7632 13024 7696 13028
rect 7712 13084 7776 13088
rect 7712 13028 7716 13084
rect 7716 13028 7772 13084
rect 7772 13028 7776 13084
rect 7712 13024 7776 13028
rect 12187 13084 12251 13088
rect 12187 13028 12191 13084
rect 12191 13028 12247 13084
rect 12247 13028 12251 13084
rect 12187 13024 12251 13028
rect 12267 13084 12331 13088
rect 12267 13028 12271 13084
rect 12271 13028 12327 13084
rect 12327 13028 12331 13084
rect 12267 13024 12331 13028
rect 12347 13084 12411 13088
rect 12347 13028 12351 13084
rect 12351 13028 12407 13084
rect 12407 13028 12411 13084
rect 12347 13024 12411 13028
rect 12427 13084 12491 13088
rect 12427 13028 12431 13084
rect 12431 13028 12487 13084
rect 12487 13028 12491 13084
rect 12427 13024 12491 13028
rect 16902 13084 16966 13088
rect 16902 13028 16906 13084
rect 16906 13028 16962 13084
rect 16962 13028 16966 13084
rect 16902 13024 16966 13028
rect 16982 13084 17046 13088
rect 16982 13028 16986 13084
rect 16986 13028 17042 13084
rect 17042 13028 17046 13084
rect 16982 13024 17046 13028
rect 17062 13084 17126 13088
rect 17062 13028 17066 13084
rect 17066 13028 17122 13084
rect 17122 13028 17126 13084
rect 17062 13024 17126 13028
rect 17142 13084 17206 13088
rect 17142 13028 17146 13084
rect 17146 13028 17202 13084
rect 17202 13028 17206 13084
rect 17142 13024 17206 13028
rect 8708 12684 8772 12748
rect 5114 12540 5178 12544
rect 5114 12484 5118 12540
rect 5118 12484 5174 12540
rect 5174 12484 5178 12540
rect 5114 12480 5178 12484
rect 5194 12540 5258 12544
rect 5194 12484 5198 12540
rect 5198 12484 5254 12540
rect 5254 12484 5258 12540
rect 5194 12480 5258 12484
rect 5274 12540 5338 12544
rect 5274 12484 5278 12540
rect 5278 12484 5334 12540
rect 5334 12484 5338 12540
rect 5274 12480 5338 12484
rect 5354 12540 5418 12544
rect 5354 12484 5358 12540
rect 5358 12484 5414 12540
rect 5414 12484 5418 12540
rect 5354 12480 5418 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 10069 12540 10133 12544
rect 10069 12484 10073 12540
rect 10073 12484 10129 12540
rect 10129 12484 10133 12540
rect 10069 12480 10133 12484
rect 14544 12540 14608 12544
rect 14544 12484 14548 12540
rect 14548 12484 14604 12540
rect 14604 12484 14608 12540
rect 14544 12480 14608 12484
rect 14624 12540 14688 12544
rect 14624 12484 14628 12540
rect 14628 12484 14684 12540
rect 14684 12484 14688 12540
rect 14624 12480 14688 12484
rect 14704 12540 14768 12544
rect 14704 12484 14708 12540
rect 14708 12484 14764 12540
rect 14764 12484 14768 12540
rect 14704 12480 14768 12484
rect 14784 12540 14848 12544
rect 14784 12484 14788 12540
rect 14788 12484 14844 12540
rect 14844 12484 14848 12540
rect 14784 12480 14848 12484
rect 19259 12540 19323 12544
rect 19259 12484 19263 12540
rect 19263 12484 19319 12540
rect 19319 12484 19323 12540
rect 19259 12480 19323 12484
rect 19339 12540 19403 12544
rect 19339 12484 19343 12540
rect 19343 12484 19399 12540
rect 19399 12484 19403 12540
rect 19339 12480 19403 12484
rect 19419 12540 19483 12544
rect 19419 12484 19423 12540
rect 19423 12484 19479 12540
rect 19479 12484 19483 12540
rect 19419 12480 19483 12484
rect 19499 12540 19563 12544
rect 19499 12484 19503 12540
rect 19503 12484 19559 12540
rect 19559 12484 19563 12540
rect 19499 12480 19563 12484
rect 2757 11996 2821 12000
rect 2757 11940 2761 11996
rect 2761 11940 2817 11996
rect 2817 11940 2821 11996
rect 2757 11936 2821 11940
rect 2837 11996 2901 12000
rect 2837 11940 2841 11996
rect 2841 11940 2897 11996
rect 2897 11940 2901 11996
rect 2837 11936 2901 11940
rect 2917 11996 2981 12000
rect 2917 11940 2921 11996
rect 2921 11940 2977 11996
rect 2977 11940 2981 11996
rect 2917 11936 2981 11940
rect 2997 11996 3061 12000
rect 2997 11940 3001 11996
rect 3001 11940 3057 11996
rect 3057 11940 3061 11996
rect 2997 11936 3061 11940
rect 7472 11996 7536 12000
rect 7472 11940 7476 11996
rect 7476 11940 7532 11996
rect 7532 11940 7536 11996
rect 7472 11936 7536 11940
rect 7552 11996 7616 12000
rect 7552 11940 7556 11996
rect 7556 11940 7612 11996
rect 7612 11940 7616 11996
rect 7552 11936 7616 11940
rect 7632 11996 7696 12000
rect 7632 11940 7636 11996
rect 7636 11940 7692 11996
rect 7692 11940 7696 11996
rect 7632 11936 7696 11940
rect 7712 11996 7776 12000
rect 7712 11940 7716 11996
rect 7716 11940 7772 11996
rect 7772 11940 7776 11996
rect 7712 11936 7776 11940
rect 12187 11996 12251 12000
rect 12187 11940 12191 11996
rect 12191 11940 12247 11996
rect 12247 11940 12251 11996
rect 12187 11936 12251 11940
rect 12267 11996 12331 12000
rect 12267 11940 12271 11996
rect 12271 11940 12327 11996
rect 12327 11940 12331 11996
rect 12267 11936 12331 11940
rect 12347 11996 12411 12000
rect 12347 11940 12351 11996
rect 12351 11940 12407 11996
rect 12407 11940 12411 11996
rect 12347 11936 12411 11940
rect 12427 11996 12491 12000
rect 12427 11940 12431 11996
rect 12431 11940 12487 11996
rect 12487 11940 12491 11996
rect 12427 11936 12491 11940
rect 16902 11996 16966 12000
rect 16902 11940 16906 11996
rect 16906 11940 16962 11996
rect 16962 11940 16966 11996
rect 16902 11936 16966 11940
rect 16982 11996 17046 12000
rect 16982 11940 16986 11996
rect 16986 11940 17042 11996
rect 17042 11940 17046 11996
rect 16982 11936 17046 11940
rect 17062 11996 17126 12000
rect 17062 11940 17066 11996
rect 17066 11940 17122 11996
rect 17122 11940 17126 11996
rect 17062 11936 17126 11940
rect 17142 11996 17206 12000
rect 17142 11940 17146 11996
rect 17146 11940 17202 11996
rect 17202 11940 17206 11996
rect 17142 11936 17206 11940
rect 17908 11732 17972 11796
rect 5114 11452 5178 11456
rect 5114 11396 5118 11452
rect 5118 11396 5174 11452
rect 5174 11396 5178 11452
rect 5114 11392 5178 11396
rect 5194 11452 5258 11456
rect 5194 11396 5198 11452
rect 5198 11396 5254 11452
rect 5254 11396 5258 11452
rect 5194 11392 5258 11396
rect 5274 11452 5338 11456
rect 5274 11396 5278 11452
rect 5278 11396 5334 11452
rect 5334 11396 5338 11452
rect 5274 11392 5338 11396
rect 5354 11452 5418 11456
rect 5354 11396 5358 11452
rect 5358 11396 5414 11452
rect 5414 11396 5418 11452
rect 5354 11392 5418 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 10069 11452 10133 11456
rect 10069 11396 10073 11452
rect 10073 11396 10129 11452
rect 10129 11396 10133 11452
rect 10069 11392 10133 11396
rect 14544 11452 14608 11456
rect 14544 11396 14548 11452
rect 14548 11396 14604 11452
rect 14604 11396 14608 11452
rect 14544 11392 14608 11396
rect 14624 11452 14688 11456
rect 14624 11396 14628 11452
rect 14628 11396 14684 11452
rect 14684 11396 14688 11452
rect 14624 11392 14688 11396
rect 14704 11452 14768 11456
rect 14704 11396 14708 11452
rect 14708 11396 14764 11452
rect 14764 11396 14768 11452
rect 14704 11392 14768 11396
rect 14784 11452 14848 11456
rect 14784 11396 14788 11452
rect 14788 11396 14844 11452
rect 14844 11396 14848 11452
rect 14784 11392 14848 11396
rect 19259 11452 19323 11456
rect 19259 11396 19263 11452
rect 19263 11396 19319 11452
rect 19319 11396 19323 11452
rect 19259 11392 19323 11396
rect 19339 11452 19403 11456
rect 19339 11396 19343 11452
rect 19343 11396 19399 11452
rect 19399 11396 19403 11452
rect 19339 11392 19403 11396
rect 19419 11452 19483 11456
rect 19419 11396 19423 11452
rect 19423 11396 19479 11452
rect 19479 11396 19483 11452
rect 19419 11392 19483 11396
rect 19499 11452 19563 11456
rect 19499 11396 19503 11452
rect 19503 11396 19559 11452
rect 19559 11396 19563 11452
rect 19499 11392 19563 11396
rect 2757 10908 2821 10912
rect 2757 10852 2761 10908
rect 2761 10852 2817 10908
rect 2817 10852 2821 10908
rect 2757 10848 2821 10852
rect 2837 10908 2901 10912
rect 2837 10852 2841 10908
rect 2841 10852 2897 10908
rect 2897 10852 2901 10908
rect 2837 10848 2901 10852
rect 2917 10908 2981 10912
rect 2917 10852 2921 10908
rect 2921 10852 2977 10908
rect 2977 10852 2981 10908
rect 2917 10848 2981 10852
rect 2997 10908 3061 10912
rect 2997 10852 3001 10908
rect 3001 10852 3057 10908
rect 3057 10852 3061 10908
rect 2997 10848 3061 10852
rect 7472 10908 7536 10912
rect 7472 10852 7476 10908
rect 7476 10852 7532 10908
rect 7532 10852 7536 10908
rect 7472 10848 7536 10852
rect 7552 10908 7616 10912
rect 7552 10852 7556 10908
rect 7556 10852 7612 10908
rect 7612 10852 7616 10908
rect 7552 10848 7616 10852
rect 7632 10908 7696 10912
rect 7632 10852 7636 10908
rect 7636 10852 7692 10908
rect 7692 10852 7696 10908
rect 7632 10848 7696 10852
rect 7712 10908 7776 10912
rect 7712 10852 7716 10908
rect 7716 10852 7772 10908
rect 7772 10852 7776 10908
rect 7712 10848 7776 10852
rect 12187 10908 12251 10912
rect 12187 10852 12191 10908
rect 12191 10852 12247 10908
rect 12247 10852 12251 10908
rect 12187 10848 12251 10852
rect 12267 10908 12331 10912
rect 12267 10852 12271 10908
rect 12271 10852 12327 10908
rect 12327 10852 12331 10908
rect 12267 10848 12331 10852
rect 12347 10908 12411 10912
rect 12347 10852 12351 10908
rect 12351 10852 12407 10908
rect 12407 10852 12411 10908
rect 12347 10848 12411 10852
rect 12427 10908 12491 10912
rect 12427 10852 12431 10908
rect 12431 10852 12487 10908
rect 12487 10852 12491 10908
rect 12427 10848 12491 10852
rect 16902 10908 16966 10912
rect 16902 10852 16906 10908
rect 16906 10852 16962 10908
rect 16962 10852 16966 10908
rect 16902 10848 16966 10852
rect 16982 10908 17046 10912
rect 16982 10852 16986 10908
rect 16986 10852 17042 10908
rect 17042 10852 17046 10908
rect 16982 10848 17046 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 5114 10364 5178 10368
rect 5114 10308 5118 10364
rect 5118 10308 5174 10364
rect 5174 10308 5178 10364
rect 5114 10304 5178 10308
rect 5194 10364 5258 10368
rect 5194 10308 5198 10364
rect 5198 10308 5254 10364
rect 5254 10308 5258 10364
rect 5194 10304 5258 10308
rect 5274 10364 5338 10368
rect 5274 10308 5278 10364
rect 5278 10308 5334 10364
rect 5334 10308 5338 10364
rect 5274 10304 5338 10308
rect 5354 10364 5418 10368
rect 5354 10308 5358 10364
rect 5358 10308 5414 10364
rect 5414 10308 5418 10364
rect 5354 10304 5418 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 10069 10364 10133 10368
rect 10069 10308 10073 10364
rect 10073 10308 10129 10364
rect 10129 10308 10133 10364
rect 10069 10304 10133 10308
rect 14544 10364 14608 10368
rect 14544 10308 14548 10364
rect 14548 10308 14604 10364
rect 14604 10308 14608 10364
rect 14544 10304 14608 10308
rect 14624 10364 14688 10368
rect 14624 10308 14628 10364
rect 14628 10308 14684 10364
rect 14684 10308 14688 10364
rect 14624 10304 14688 10308
rect 14704 10364 14768 10368
rect 14704 10308 14708 10364
rect 14708 10308 14764 10364
rect 14764 10308 14768 10364
rect 14704 10304 14768 10308
rect 14784 10364 14848 10368
rect 14784 10308 14788 10364
rect 14788 10308 14844 10364
rect 14844 10308 14848 10364
rect 14784 10304 14848 10308
rect 19259 10364 19323 10368
rect 19259 10308 19263 10364
rect 19263 10308 19319 10364
rect 19319 10308 19323 10364
rect 19259 10304 19323 10308
rect 19339 10364 19403 10368
rect 19339 10308 19343 10364
rect 19343 10308 19399 10364
rect 19399 10308 19403 10364
rect 19339 10304 19403 10308
rect 19419 10364 19483 10368
rect 19419 10308 19423 10364
rect 19423 10308 19479 10364
rect 19479 10308 19483 10364
rect 19419 10304 19483 10308
rect 19499 10364 19563 10368
rect 19499 10308 19503 10364
rect 19503 10308 19559 10364
rect 19559 10308 19563 10364
rect 19499 10304 19563 10308
rect 2757 9820 2821 9824
rect 2757 9764 2761 9820
rect 2761 9764 2817 9820
rect 2817 9764 2821 9820
rect 2757 9760 2821 9764
rect 2837 9820 2901 9824
rect 2837 9764 2841 9820
rect 2841 9764 2897 9820
rect 2897 9764 2901 9820
rect 2837 9760 2901 9764
rect 2917 9820 2981 9824
rect 2917 9764 2921 9820
rect 2921 9764 2977 9820
rect 2977 9764 2981 9820
rect 2917 9760 2981 9764
rect 2997 9820 3061 9824
rect 2997 9764 3001 9820
rect 3001 9764 3057 9820
rect 3057 9764 3061 9820
rect 2997 9760 3061 9764
rect 7472 9820 7536 9824
rect 7472 9764 7476 9820
rect 7476 9764 7532 9820
rect 7532 9764 7536 9820
rect 7472 9760 7536 9764
rect 7552 9820 7616 9824
rect 7552 9764 7556 9820
rect 7556 9764 7612 9820
rect 7612 9764 7616 9820
rect 7552 9760 7616 9764
rect 7632 9820 7696 9824
rect 7632 9764 7636 9820
rect 7636 9764 7692 9820
rect 7692 9764 7696 9820
rect 7632 9760 7696 9764
rect 7712 9820 7776 9824
rect 7712 9764 7716 9820
rect 7716 9764 7772 9820
rect 7772 9764 7776 9820
rect 7712 9760 7776 9764
rect 12187 9820 12251 9824
rect 12187 9764 12191 9820
rect 12191 9764 12247 9820
rect 12247 9764 12251 9820
rect 12187 9760 12251 9764
rect 12267 9820 12331 9824
rect 12267 9764 12271 9820
rect 12271 9764 12327 9820
rect 12327 9764 12331 9820
rect 12267 9760 12331 9764
rect 12347 9820 12411 9824
rect 12347 9764 12351 9820
rect 12351 9764 12407 9820
rect 12407 9764 12411 9820
rect 12347 9760 12411 9764
rect 12427 9820 12491 9824
rect 12427 9764 12431 9820
rect 12431 9764 12487 9820
rect 12487 9764 12491 9820
rect 12427 9760 12491 9764
rect 16902 9820 16966 9824
rect 16902 9764 16906 9820
rect 16906 9764 16962 9820
rect 16962 9764 16966 9820
rect 16902 9760 16966 9764
rect 16982 9820 17046 9824
rect 16982 9764 16986 9820
rect 16986 9764 17042 9820
rect 17042 9764 17046 9820
rect 16982 9760 17046 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 5114 9276 5178 9280
rect 5114 9220 5118 9276
rect 5118 9220 5174 9276
rect 5174 9220 5178 9276
rect 5114 9216 5178 9220
rect 5194 9276 5258 9280
rect 5194 9220 5198 9276
rect 5198 9220 5254 9276
rect 5254 9220 5258 9276
rect 5194 9216 5258 9220
rect 5274 9276 5338 9280
rect 5274 9220 5278 9276
rect 5278 9220 5334 9276
rect 5334 9220 5338 9276
rect 5274 9216 5338 9220
rect 5354 9276 5418 9280
rect 5354 9220 5358 9276
rect 5358 9220 5414 9276
rect 5414 9220 5418 9276
rect 5354 9216 5418 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 10069 9276 10133 9280
rect 10069 9220 10073 9276
rect 10073 9220 10129 9276
rect 10129 9220 10133 9276
rect 10069 9216 10133 9220
rect 14544 9276 14608 9280
rect 14544 9220 14548 9276
rect 14548 9220 14604 9276
rect 14604 9220 14608 9276
rect 14544 9216 14608 9220
rect 14624 9276 14688 9280
rect 14624 9220 14628 9276
rect 14628 9220 14684 9276
rect 14684 9220 14688 9276
rect 14624 9216 14688 9220
rect 14704 9276 14768 9280
rect 14704 9220 14708 9276
rect 14708 9220 14764 9276
rect 14764 9220 14768 9276
rect 14704 9216 14768 9220
rect 14784 9276 14848 9280
rect 14784 9220 14788 9276
rect 14788 9220 14844 9276
rect 14844 9220 14848 9276
rect 14784 9216 14848 9220
rect 19259 9276 19323 9280
rect 19259 9220 19263 9276
rect 19263 9220 19319 9276
rect 19319 9220 19323 9276
rect 19259 9216 19323 9220
rect 19339 9276 19403 9280
rect 19339 9220 19343 9276
rect 19343 9220 19399 9276
rect 19399 9220 19403 9276
rect 19339 9216 19403 9220
rect 19419 9276 19483 9280
rect 19419 9220 19423 9276
rect 19423 9220 19479 9276
rect 19479 9220 19483 9276
rect 19419 9216 19483 9220
rect 19499 9276 19563 9280
rect 19499 9220 19503 9276
rect 19503 9220 19559 9276
rect 19559 9220 19563 9276
rect 19499 9216 19563 9220
rect 2757 8732 2821 8736
rect 2757 8676 2761 8732
rect 2761 8676 2817 8732
rect 2817 8676 2821 8732
rect 2757 8672 2821 8676
rect 2837 8732 2901 8736
rect 2837 8676 2841 8732
rect 2841 8676 2897 8732
rect 2897 8676 2901 8732
rect 2837 8672 2901 8676
rect 2917 8732 2981 8736
rect 2917 8676 2921 8732
rect 2921 8676 2977 8732
rect 2977 8676 2981 8732
rect 2917 8672 2981 8676
rect 2997 8732 3061 8736
rect 2997 8676 3001 8732
rect 3001 8676 3057 8732
rect 3057 8676 3061 8732
rect 2997 8672 3061 8676
rect 7472 8732 7536 8736
rect 7472 8676 7476 8732
rect 7476 8676 7532 8732
rect 7532 8676 7536 8732
rect 7472 8672 7536 8676
rect 7552 8732 7616 8736
rect 7552 8676 7556 8732
rect 7556 8676 7612 8732
rect 7612 8676 7616 8732
rect 7552 8672 7616 8676
rect 7632 8732 7696 8736
rect 7632 8676 7636 8732
rect 7636 8676 7692 8732
rect 7692 8676 7696 8732
rect 7632 8672 7696 8676
rect 7712 8732 7776 8736
rect 7712 8676 7716 8732
rect 7716 8676 7772 8732
rect 7772 8676 7776 8732
rect 7712 8672 7776 8676
rect 12187 8732 12251 8736
rect 12187 8676 12191 8732
rect 12191 8676 12247 8732
rect 12247 8676 12251 8732
rect 12187 8672 12251 8676
rect 12267 8732 12331 8736
rect 12267 8676 12271 8732
rect 12271 8676 12327 8732
rect 12327 8676 12331 8732
rect 12267 8672 12331 8676
rect 12347 8732 12411 8736
rect 12347 8676 12351 8732
rect 12351 8676 12407 8732
rect 12407 8676 12411 8732
rect 12347 8672 12411 8676
rect 12427 8732 12491 8736
rect 12427 8676 12431 8732
rect 12431 8676 12487 8732
rect 12487 8676 12491 8732
rect 12427 8672 12491 8676
rect 16902 8732 16966 8736
rect 16902 8676 16906 8732
rect 16906 8676 16962 8732
rect 16962 8676 16966 8732
rect 16902 8672 16966 8676
rect 16982 8732 17046 8736
rect 16982 8676 16986 8732
rect 16986 8676 17042 8732
rect 17042 8676 17046 8732
rect 16982 8672 17046 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 5114 8188 5178 8192
rect 5114 8132 5118 8188
rect 5118 8132 5174 8188
rect 5174 8132 5178 8188
rect 5114 8128 5178 8132
rect 5194 8188 5258 8192
rect 5194 8132 5198 8188
rect 5198 8132 5254 8188
rect 5254 8132 5258 8188
rect 5194 8128 5258 8132
rect 5274 8188 5338 8192
rect 5274 8132 5278 8188
rect 5278 8132 5334 8188
rect 5334 8132 5338 8188
rect 5274 8128 5338 8132
rect 5354 8188 5418 8192
rect 5354 8132 5358 8188
rect 5358 8132 5414 8188
rect 5414 8132 5418 8188
rect 5354 8128 5418 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 10069 8188 10133 8192
rect 10069 8132 10073 8188
rect 10073 8132 10129 8188
rect 10129 8132 10133 8188
rect 10069 8128 10133 8132
rect 14544 8188 14608 8192
rect 14544 8132 14548 8188
rect 14548 8132 14604 8188
rect 14604 8132 14608 8188
rect 14544 8128 14608 8132
rect 14624 8188 14688 8192
rect 14624 8132 14628 8188
rect 14628 8132 14684 8188
rect 14684 8132 14688 8188
rect 14624 8128 14688 8132
rect 14704 8188 14768 8192
rect 14704 8132 14708 8188
rect 14708 8132 14764 8188
rect 14764 8132 14768 8188
rect 14704 8128 14768 8132
rect 14784 8188 14848 8192
rect 14784 8132 14788 8188
rect 14788 8132 14844 8188
rect 14844 8132 14848 8188
rect 14784 8128 14848 8132
rect 19259 8188 19323 8192
rect 19259 8132 19263 8188
rect 19263 8132 19319 8188
rect 19319 8132 19323 8188
rect 19259 8128 19323 8132
rect 19339 8188 19403 8192
rect 19339 8132 19343 8188
rect 19343 8132 19399 8188
rect 19399 8132 19403 8188
rect 19339 8128 19403 8132
rect 19419 8188 19483 8192
rect 19419 8132 19423 8188
rect 19423 8132 19479 8188
rect 19479 8132 19483 8188
rect 19419 8128 19483 8132
rect 19499 8188 19563 8192
rect 19499 8132 19503 8188
rect 19503 8132 19559 8188
rect 19559 8132 19563 8188
rect 19499 8128 19563 8132
rect 2757 7644 2821 7648
rect 2757 7588 2761 7644
rect 2761 7588 2817 7644
rect 2817 7588 2821 7644
rect 2757 7584 2821 7588
rect 2837 7644 2901 7648
rect 2837 7588 2841 7644
rect 2841 7588 2897 7644
rect 2897 7588 2901 7644
rect 2837 7584 2901 7588
rect 2917 7644 2981 7648
rect 2917 7588 2921 7644
rect 2921 7588 2977 7644
rect 2977 7588 2981 7644
rect 2917 7584 2981 7588
rect 2997 7644 3061 7648
rect 2997 7588 3001 7644
rect 3001 7588 3057 7644
rect 3057 7588 3061 7644
rect 2997 7584 3061 7588
rect 7472 7644 7536 7648
rect 7472 7588 7476 7644
rect 7476 7588 7532 7644
rect 7532 7588 7536 7644
rect 7472 7584 7536 7588
rect 7552 7644 7616 7648
rect 7552 7588 7556 7644
rect 7556 7588 7612 7644
rect 7612 7588 7616 7644
rect 7552 7584 7616 7588
rect 7632 7644 7696 7648
rect 7632 7588 7636 7644
rect 7636 7588 7692 7644
rect 7692 7588 7696 7644
rect 7632 7584 7696 7588
rect 7712 7644 7776 7648
rect 7712 7588 7716 7644
rect 7716 7588 7772 7644
rect 7772 7588 7776 7644
rect 7712 7584 7776 7588
rect 12187 7644 12251 7648
rect 12187 7588 12191 7644
rect 12191 7588 12247 7644
rect 12247 7588 12251 7644
rect 12187 7584 12251 7588
rect 12267 7644 12331 7648
rect 12267 7588 12271 7644
rect 12271 7588 12327 7644
rect 12327 7588 12331 7644
rect 12267 7584 12331 7588
rect 12347 7644 12411 7648
rect 12347 7588 12351 7644
rect 12351 7588 12407 7644
rect 12407 7588 12411 7644
rect 12347 7584 12411 7588
rect 12427 7644 12491 7648
rect 12427 7588 12431 7644
rect 12431 7588 12487 7644
rect 12487 7588 12491 7644
rect 12427 7584 12491 7588
rect 16902 7644 16966 7648
rect 16902 7588 16906 7644
rect 16906 7588 16962 7644
rect 16962 7588 16966 7644
rect 16902 7584 16966 7588
rect 16982 7644 17046 7648
rect 16982 7588 16986 7644
rect 16986 7588 17042 7644
rect 17042 7588 17046 7644
rect 16982 7584 17046 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 5114 7100 5178 7104
rect 5114 7044 5118 7100
rect 5118 7044 5174 7100
rect 5174 7044 5178 7100
rect 5114 7040 5178 7044
rect 5194 7100 5258 7104
rect 5194 7044 5198 7100
rect 5198 7044 5254 7100
rect 5254 7044 5258 7100
rect 5194 7040 5258 7044
rect 5274 7100 5338 7104
rect 5274 7044 5278 7100
rect 5278 7044 5334 7100
rect 5334 7044 5338 7100
rect 5274 7040 5338 7044
rect 5354 7100 5418 7104
rect 5354 7044 5358 7100
rect 5358 7044 5414 7100
rect 5414 7044 5418 7100
rect 5354 7040 5418 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 10069 7100 10133 7104
rect 10069 7044 10073 7100
rect 10073 7044 10129 7100
rect 10129 7044 10133 7100
rect 10069 7040 10133 7044
rect 14544 7100 14608 7104
rect 14544 7044 14548 7100
rect 14548 7044 14604 7100
rect 14604 7044 14608 7100
rect 14544 7040 14608 7044
rect 14624 7100 14688 7104
rect 14624 7044 14628 7100
rect 14628 7044 14684 7100
rect 14684 7044 14688 7100
rect 14624 7040 14688 7044
rect 14704 7100 14768 7104
rect 14704 7044 14708 7100
rect 14708 7044 14764 7100
rect 14764 7044 14768 7100
rect 14704 7040 14768 7044
rect 14784 7100 14848 7104
rect 14784 7044 14788 7100
rect 14788 7044 14844 7100
rect 14844 7044 14848 7100
rect 14784 7040 14848 7044
rect 19259 7100 19323 7104
rect 19259 7044 19263 7100
rect 19263 7044 19319 7100
rect 19319 7044 19323 7100
rect 19259 7040 19323 7044
rect 19339 7100 19403 7104
rect 19339 7044 19343 7100
rect 19343 7044 19399 7100
rect 19399 7044 19403 7100
rect 19339 7040 19403 7044
rect 19419 7100 19483 7104
rect 19419 7044 19423 7100
rect 19423 7044 19479 7100
rect 19479 7044 19483 7100
rect 19419 7040 19483 7044
rect 19499 7100 19563 7104
rect 19499 7044 19503 7100
rect 19503 7044 19559 7100
rect 19559 7044 19563 7100
rect 19499 7040 19563 7044
rect 10364 6836 10428 6900
rect 2757 6556 2821 6560
rect 2757 6500 2761 6556
rect 2761 6500 2817 6556
rect 2817 6500 2821 6556
rect 2757 6496 2821 6500
rect 2837 6556 2901 6560
rect 2837 6500 2841 6556
rect 2841 6500 2897 6556
rect 2897 6500 2901 6556
rect 2837 6496 2901 6500
rect 2917 6556 2981 6560
rect 2917 6500 2921 6556
rect 2921 6500 2977 6556
rect 2977 6500 2981 6556
rect 2917 6496 2981 6500
rect 2997 6556 3061 6560
rect 2997 6500 3001 6556
rect 3001 6500 3057 6556
rect 3057 6500 3061 6556
rect 2997 6496 3061 6500
rect 7472 6556 7536 6560
rect 7472 6500 7476 6556
rect 7476 6500 7532 6556
rect 7532 6500 7536 6556
rect 7472 6496 7536 6500
rect 7552 6556 7616 6560
rect 7552 6500 7556 6556
rect 7556 6500 7612 6556
rect 7612 6500 7616 6556
rect 7552 6496 7616 6500
rect 7632 6556 7696 6560
rect 7632 6500 7636 6556
rect 7636 6500 7692 6556
rect 7692 6500 7696 6556
rect 7632 6496 7696 6500
rect 7712 6556 7776 6560
rect 7712 6500 7716 6556
rect 7716 6500 7772 6556
rect 7772 6500 7776 6556
rect 7712 6496 7776 6500
rect 12187 6556 12251 6560
rect 12187 6500 12191 6556
rect 12191 6500 12247 6556
rect 12247 6500 12251 6556
rect 12187 6496 12251 6500
rect 12267 6556 12331 6560
rect 12267 6500 12271 6556
rect 12271 6500 12327 6556
rect 12327 6500 12331 6556
rect 12267 6496 12331 6500
rect 12347 6556 12411 6560
rect 12347 6500 12351 6556
rect 12351 6500 12407 6556
rect 12407 6500 12411 6556
rect 12347 6496 12411 6500
rect 12427 6556 12491 6560
rect 12427 6500 12431 6556
rect 12431 6500 12487 6556
rect 12487 6500 12491 6556
rect 12427 6496 12491 6500
rect 16902 6556 16966 6560
rect 16902 6500 16906 6556
rect 16906 6500 16962 6556
rect 16962 6500 16966 6556
rect 16902 6496 16966 6500
rect 16982 6556 17046 6560
rect 16982 6500 16986 6556
rect 16986 6500 17042 6556
rect 17042 6500 17046 6556
rect 16982 6496 17046 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 5114 6012 5178 6016
rect 5114 5956 5118 6012
rect 5118 5956 5174 6012
rect 5174 5956 5178 6012
rect 5114 5952 5178 5956
rect 5194 6012 5258 6016
rect 5194 5956 5198 6012
rect 5198 5956 5254 6012
rect 5254 5956 5258 6012
rect 5194 5952 5258 5956
rect 5274 6012 5338 6016
rect 5274 5956 5278 6012
rect 5278 5956 5334 6012
rect 5334 5956 5338 6012
rect 5274 5952 5338 5956
rect 5354 6012 5418 6016
rect 5354 5956 5358 6012
rect 5358 5956 5414 6012
rect 5414 5956 5418 6012
rect 5354 5952 5418 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 10069 6012 10133 6016
rect 10069 5956 10073 6012
rect 10073 5956 10129 6012
rect 10129 5956 10133 6012
rect 10069 5952 10133 5956
rect 14544 6012 14608 6016
rect 14544 5956 14548 6012
rect 14548 5956 14604 6012
rect 14604 5956 14608 6012
rect 14544 5952 14608 5956
rect 14624 6012 14688 6016
rect 14624 5956 14628 6012
rect 14628 5956 14684 6012
rect 14684 5956 14688 6012
rect 14624 5952 14688 5956
rect 14704 6012 14768 6016
rect 14704 5956 14708 6012
rect 14708 5956 14764 6012
rect 14764 5956 14768 6012
rect 14704 5952 14768 5956
rect 14784 6012 14848 6016
rect 14784 5956 14788 6012
rect 14788 5956 14844 6012
rect 14844 5956 14848 6012
rect 14784 5952 14848 5956
rect 19259 6012 19323 6016
rect 19259 5956 19263 6012
rect 19263 5956 19319 6012
rect 19319 5956 19323 6012
rect 19259 5952 19323 5956
rect 19339 6012 19403 6016
rect 19339 5956 19343 6012
rect 19343 5956 19399 6012
rect 19399 5956 19403 6012
rect 19339 5952 19403 5956
rect 19419 6012 19483 6016
rect 19419 5956 19423 6012
rect 19423 5956 19479 6012
rect 19479 5956 19483 6012
rect 19419 5952 19483 5956
rect 19499 6012 19563 6016
rect 19499 5956 19503 6012
rect 19503 5956 19559 6012
rect 19559 5956 19563 6012
rect 19499 5952 19563 5956
rect 2757 5468 2821 5472
rect 2757 5412 2761 5468
rect 2761 5412 2817 5468
rect 2817 5412 2821 5468
rect 2757 5408 2821 5412
rect 2837 5468 2901 5472
rect 2837 5412 2841 5468
rect 2841 5412 2897 5468
rect 2897 5412 2901 5468
rect 2837 5408 2901 5412
rect 2917 5468 2981 5472
rect 2917 5412 2921 5468
rect 2921 5412 2977 5468
rect 2977 5412 2981 5468
rect 2917 5408 2981 5412
rect 2997 5468 3061 5472
rect 2997 5412 3001 5468
rect 3001 5412 3057 5468
rect 3057 5412 3061 5468
rect 2997 5408 3061 5412
rect 7472 5468 7536 5472
rect 7472 5412 7476 5468
rect 7476 5412 7532 5468
rect 7532 5412 7536 5468
rect 7472 5408 7536 5412
rect 7552 5468 7616 5472
rect 7552 5412 7556 5468
rect 7556 5412 7612 5468
rect 7612 5412 7616 5468
rect 7552 5408 7616 5412
rect 7632 5468 7696 5472
rect 7632 5412 7636 5468
rect 7636 5412 7692 5468
rect 7692 5412 7696 5468
rect 7632 5408 7696 5412
rect 7712 5468 7776 5472
rect 7712 5412 7716 5468
rect 7716 5412 7772 5468
rect 7772 5412 7776 5468
rect 7712 5408 7776 5412
rect 12187 5468 12251 5472
rect 12187 5412 12191 5468
rect 12191 5412 12247 5468
rect 12247 5412 12251 5468
rect 12187 5408 12251 5412
rect 12267 5468 12331 5472
rect 12267 5412 12271 5468
rect 12271 5412 12327 5468
rect 12327 5412 12331 5468
rect 12267 5408 12331 5412
rect 12347 5468 12411 5472
rect 12347 5412 12351 5468
rect 12351 5412 12407 5468
rect 12407 5412 12411 5468
rect 12347 5408 12411 5412
rect 12427 5468 12491 5472
rect 12427 5412 12431 5468
rect 12431 5412 12487 5468
rect 12487 5412 12491 5468
rect 12427 5408 12491 5412
rect 16902 5468 16966 5472
rect 16902 5412 16906 5468
rect 16906 5412 16962 5468
rect 16962 5412 16966 5468
rect 16902 5408 16966 5412
rect 16982 5468 17046 5472
rect 16982 5412 16986 5468
rect 16986 5412 17042 5468
rect 17042 5412 17046 5468
rect 16982 5408 17046 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 5114 4924 5178 4928
rect 5114 4868 5118 4924
rect 5118 4868 5174 4924
rect 5174 4868 5178 4924
rect 5114 4864 5178 4868
rect 5194 4924 5258 4928
rect 5194 4868 5198 4924
rect 5198 4868 5254 4924
rect 5254 4868 5258 4924
rect 5194 4864 5258 4868
rect 5274 4924 5338 4928
rect 5274 4868 5278 4924
rect 5278 4868 5334 4924
rect 5334 4868 5338 4924
rect 5274 4864 5338 4868
rect 5354 4924 5418 4928
rect 5354 4868 5358 4924
rect 5358 4868 5414 4924
rect 5414 4868 5418 4924
rect 5354 4864 5418 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 10069 4924 10133 4928
rect 10069 4868 10073 4924
rect 10073 4868 10129 4924
rect 10129 4868 10133 4924
rect 10069 4864 10133 4868
rect 14544 4924 14608 4928
rect 14544 4868 14548 4924
rect 14548 4868 14604 4924
rect 14604 4868 14608 4924
rect 14544 4864 14608 4868
rect 14624 4924 14688 4928
rect 14624 4868 14628 4924
rect 14628 4868 14684 4924
rect 14684 4868 14688 4924
rect 14624 4864 14688 4868
rect 14704 4924 14768 4928
rect 14704 4868 14708 4924
rect 14708 4868 14764 4924
rect 14764 4868 14768 4924
rect 14704 4864 14768 4868
rect 14784 4924 14848 4928
rect 14784 4868 14788 4924
rect 14788 4868 14844 4924
rect 14844 4868 14848 4924
rect 14784 4864 14848 4868
rect 19259 4924 19323 4928
rect 19259 4868 19263 4924
rect 19263 4868 19319 4924
rect 19319 4868 19323 4924
rect 19259 4864 19323 4868
rect 19339 4924 19403 4928
rect 19339 4868 19343 4924
rect 19343 4868 19399 4924
rect 19399 4868 19403 4924
rect 19339 4864 19403 4868
rect 19419 4924 19483 4928
rect 19419 4868 19423 4924
rect 19423 4868 19479 4924
rect 19479 4868 19483 4924
rect 19419 4864 19483 4868
rect 19499 4924 19563 4928
rect 19499 4868 19503 4924
rect 19503 4868 19559 4924
rect 19559 4868 19563 4924
rect 19499 4864 19563 4868
rect 2757 4380 2821 4384
rect 2757 4324 2761 4380
rect 2761 4324 2817 4380
rect 2817 4324 2821 4380
rect 2757 4320 2821 4324
rect 2837 4380 2901 4384
rect 2837 4324 2841 4380
rect 2841 4324 2897 4380
rect 2897 4324 2901 4380
rect 2837 4320 2901 4324
rect 2917 4380 2981 4384
rect 2917 4324 2921 4380
rect 2921 4324 2977 4380
rect 2977 4324 2981 4380
rect 2917 4320 2981 4324
rect 2997 4380 3061 4384
rect 2997 4324 3001 4380
rect 3001 4324 3057 4380
rect 3057 4324 3061 4380
rect 2997 4320 3061 4324
rect 7472 4380 7536 4384
rect 7472 4324 7476 4380
rect 7476 4324 7532 4380
rect 7532 4324 7536 4380
rect 7472 4320 7536 4324
rect 7552 4380 7616 4384
rect 7552 4324 7556 4380
rect 7556 4324 7612 4380
rect 7612 4324 7616 4380
rect 7552 4320 7616 4324
rect 7632 4380 7696 4384
rect 7632 4324 7636 4380
rect 7636 4324 7692 4380
rect 7692 4324 7696 4380
rect 7632 4320 7696 4324
rect 7712 4380 7776 4384
rect 7712 4324 7716 4380
rect 7716 4324 7772 4380
rect 7772 4324 7776 4380
rect 7712 4320 7776 4324
rect 12187 4380 12251 4384
rect 12187 4324 12191 4380
rect 12191 4324 12247 4380
rect 12247 4324 12251 4380
rect 12187 4320 12251 4324
rect 12267 4380 12331 4384
rect 12267 4324 12271 4380
rect 12271 4324 12327 4380
rect 12327 4324 12331 4380
rect 12267 4320 12331 4324
rect 12347 4380 12411 4384
rect 12347 4324 12351 4380
rect 12351 4324 12407 4380
rect 12407 4324 12411 4380
rect 12347 4320 12411 4324
rect 12427 4380 12491 4384
rect 12427 4324 12431 4380
rect 12431 4324 12487 4380
rect 12487 4324 12491 4380
rect 12427 4320 12491 4324
rect 16902 4380 16966 4384
rect 16902 4324 16906 4380
rect 16906 4324 16962 4380
rect 16962 4324 16966 4380
rect 16902 4320 16966 4324
rect 16982 4380 17046 4384
rect 16982 4324 16986 4380
rect 16986 4324 17042 4380
rect 17042 4324 17046 4380
rect 16982 4320 17046 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 5114 3836 5178 3840
rect 5114 3780 5118 3836
rect 5118 3780 5174 3836
rect 5174 3780 5178 3836
rect 5114 3776 5178 3780
rect 5194 3836 5258 3840
rect 5194 3780 5198 3836
rect 5198 3780 5254 3836
rect 5254 3780 5258 3836
rect 5194 3776 5258 3780
rect 5274 3836 5338 3840
rect 5274 3780 5278 3836
rect 5278 3780 5334 3836
rect 5334 3780 5338 3836
rect 5274 3776 5338 3780
rect 5354 3836 5418 3840
rect 5354 3780 5358 3836
rect 5358 3780 5414 3836
rect 5414 3780 5418 3836
rect 5354 3776 5418 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 10069 3836 10133 3840
rect 10069 3780 10073 3836
rect 10073 3780 10129 3836
rect 10129 3780 10133 3836
rect 10069 3776 10133 3780
rect 14544 3836 14608 3840
rect 14544 3780 14548 3836
rect 14548 3780 14604 3836
rect 14604 3780 14608 3836
rect 14544 3776 14608 3780
rect 14624 3836 14688 3840
rect 14624 3780 14628 3836
rect 14628 3780 14684 3836
rect 14684 3780 14688 3836
rect 14624 3776 14688 3780
rect 14704 3836 14768 3840
rect 14704 3780 14708 3836
rect 14708 3780 14764 3836
rect 14764 3780 14768 3836
rect 14704 3776 14768 3780
rect 14784 3836 14848 3840
rect 14784 3780 14788 3836
rect 14788 3780 14844 3836
rect 14844 3780 14848 3836
rect 14784 3776 14848 3780
rect 19259 3836 19323 3840
rect 19259 3780 19263 3836
rect 19263 3780 19319 3836
rect 19319 3780 19323 3836
rect 19259 3776 19323 3780
rect 19339 3836 19403 3840
rect 19339 3780 19343 3836
rect 19343 3780 19399 3836
rect 19399 3780 19403 3836
rect 19339 3776 19403 3780
rect 19419 3836 19483 3840
rect 19419 3780 19423 3836
rect 19423 3780 19479 3836
rect 19479 3780 19483 3836
rect 19419 3776 19483 3780
rect 19499 3836 19563 3840
rect 19499 3780 19503 3836
rect 19503 3780 19559 3836
rect 19559 3780 19563 3836
rect 19499 3776 19563 3780
rect 2757 3292 2821 3296
rect 2757 3236 2761 3292
rect 2761 3236 2817 3292
rect 2817 3236 2821 3292
rect 2757 3232 2821 3236
rect 2837 3292 2901 3296
rect 2837 3236 2841 3292
rect 2841 3236 2897 3292
rect 2897 3236 2901 3292
rect 2837 3232 2901 3236
rect 2917 3292 2981 3296
rect 2917 3236 2921 3292
rect 2921 3236 2977 3292
rect 2977 3236 2981 3292
rect 2917 3232 2981 3236
rect 2997 3292 3061 3296
rect 2997 3236 3001 3292
rect 3001 3236 3057 3292
rect 3057 3236 3061 3292
rect 2997 3232 3061 3236
rect 7472 3292 7536 3296
rect 7472 3236 7476 3292
rect 7476 3236 7532 3292
rect 7532 3236 7536 3292
rect 7472 3232 7536 3236
rect 7552 3292 7616 3296
rect 7552 3236 7556 3292
rect 7556 3236 7612 3292
rect 7612 3236 7616 3292
rect 7552 3232 7616 3236
rect 7632 3292 7696 3296
rect 7632 3236 7636 3292
rect 7636 3236 7692 3292
rect 7692 3236 7696 3292
rect 7632 3232 7696 3236
rect 7712 3292 7776 3296
rect 7712 3236 7716 3292
rect 7716 3236 7772 3292
rect 7772 3236 7776 3292
rect 7712 3232 7776 3236
rect 12187 3292 12251 3296
rect 12187 3236 12191 3292
rect 12191 3236 12247 3292
rect 12247 3236 12251 3292
rect 12187 3232 12251 3236
rect 12267 3292 12331 3296
rect 12267 3236 12271 3292
rect 12271 3236 12327 3292
rect 12327 3236 12331 3292
rect 12267 3232 12331 3236
rect 12347 3292 12411 3296
rect 12347 3236 12351 3292
rect 12351 3236 12407 3292
rect 12407 3236 12411 3292
rect 12347 3232 12411 3236
rect 12427 3292 12491 3296
rect 12427 3236 12431 3292
rect 12431 3236 12487 3292
rect 12487 3236 12491 3292
rect 12427 3232 12491 3236
rect 16902 3292 16966 3296
rect 16902 3236 16906 3292
rect 16906 3236 16962 3292
rect 16962 3236 16966 3292
rect 16902 3232 16966 3236
rect 16982 3292 17046 3296
rect 16982 3236 16986 3292
rect 16986 3236 17042 3292
rect 17042 3236 17046 3292
rect 16982 3232 17046 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 5114 2748 5178 2752
rect 5114 2692 5118 2748
rect 5118 2692 5174 2748
rect 5174 2692 5178 2748
rect 5114 2688 5178 2692
rect 5194 2748 5258 2752
rect 5194 2692 5198 2748
rect 5198 2692 5254 2748
rect 5254 2692 5258 2748
rect 5194 2688 5258 2692
rect 5274 2748 5338 2752
rect 5274 2692 5278 2748
rect 5278 2692 5334 2748
rect 5334 2692 5338 2748
rect 5274 2688 5338 2692
rect 5354 2748 5418 2752
rect 5354 2692 5358 2748
rect 5358 2692 5414 2748
rect 5414 2692 5418 2748
rect 5354 2688 5418 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 10069 2748 10133 2752
rect 10069 2692 10073 2748
rect 10073 2692 10129 2748
rect 10129 2692 10133 2748
rect 10069 2688 10133 2692
rect 14544 2748 14608 2752
rect 14544 2692 14548 2748
rect 14548 2692 14604 2748
rect 14604 2692 14608 2748
rect 14544 2688 14608 2692
rect 14624 2748 14688 2752
rect 14624 2692 14628 2748
rect 14628 2692 14684 2748
rect 14684 2692 14688 2748
rect 14624 2688 14688 2692
rect 14704 2748 14768 2752
rect 14704 2692 14708 2748
rect 14708 2692 14764 2748
rect 14764 2692 14768 2748
rect 14704 2688 14768 2692
rect 14784 2748 14848 2752
rect 14784 2692 14788 2748
rect 14788 2692 14844 2748
rect 14844 2692 14848 2748
rect 14784 2688 14848 2692
rect 19259 2748 19323 2752
rect 19259 2692 19263 2748
rect 19263 2692 19319 2748
rect 19319 2692 19323 2748
rect 19259 2688 19323 2692
rect 19339 2748 19403 2752
rect 19339 2692 19343 2748
rect 19343 2692 19399 2748
rect 19399 2692 19403 2748
rect 19339 2688 19403 2692
rect 19419 2748 19483 2752
rect 19419 2692 19423 2748
rect 19423 2692 19479 2748
rect 19479 2692 19483 2748
rect 19419 2688 19483 2692
rect 19499 2748 19563 2752
rect 19499 2692 19503 2748
rect 19503 2692 19559 2748
rect 19559 2692 19563 2748
rect 19499 2688 19563 2692
rect 2757 2204 2821 2208
rect 2757 2148 2761 2204
rect 2761 2148 2817 2204
rect 2817 2148 2821 2204
rect 2757 2144 2821 2148
rect 2837 2204 2901 2208
rect 2837 2148 2841 2204
rect 2841 2148 2897 2204
rect 2897 2148 2901 2204
rect 2837 2144 2901 2148
rect 2917 2204 2981 2208
rect 2917 2148 2921 2204
rect 2921 2148 2977 2204
rect 2977 2148 2981 2204
rect 2917 2144 2981 2148
rect 2997 2204 3061 2208
rect 2997 2148 3001 2204
rect 3001 2148 3057 2204
rect 3057 2148 3061 2204
rect 2997 2144 3061 2148
rect 7472 2204 7536 2208
rect 7472 2148 7476 2204
rect 7476 2148 7532 2204
rect 7532 2148 7536 2204
rect 7472 2144 7536 2148
rect 7552 2204 7616 2208
rect 7552 2148 7556 2204
rect 7556 2148 7612 2204
rect 7612 2148 7616 2204
rect 7552 2144 7616 2148
rect 7632 2204 7696 2208
rect 7632 2148 7636 2204
rect 7636 2148 7692 2204
rect 7692 2148 7696 2204
rect 7632 2144 7696 2148
rect 7712 2204 7776 2208
rect 7712 2148 7716 2204
rect 7716 2148 7772 2204
rect 7772 2148 7776 2204
rect 7712 2144 7776 2148
rect 12187 2204 12251 2208
rect 12187 2148 12191 2204
rect 12191 2148 12247 2204
rect 12247 2148 12251 2204
rect 12187 2144 12251 2148
rect 12267 2204 12331 2208
rect 12267 2148 12271 2204
rect 12271 2148 12327 2204
rect 12327 2148 12331 2204
rect 12267 2144 12331 2148
rect 12347 2204 12411 2208
rect 12347 2148 12351 2204
rect 12351 2148 12407 2204
rect 12407 2148 12411 2204
rect 12347 2144 12411 2148
rect 12427 2204 12491 2208
rect 12427 2148 12431 2204
rect 12431 2148 12487 2204
rect 12487 2148 12491 2204
rect 12427 2144 12491 2148
rect 16902 2204 16966 2208
rect 16902 2148 16906 2204
rect 16906 2148 16962 2204
rect 16962 2148 16966 2204
rect 16902 2144 16966 2148
rect 16982 2204 17046 2208
rect 16982 2148 16986 2204
rect 16986 2148 17042 2204
rect 17042 2148 17046 2204
rect 16982 2144 17046 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 5114 1660 5178 1664
rect 5114 1604 5118 1660
rect 5118 1604 5174 1660
rect 5174 1604 5178 1660
rect 5114 1600 5178 1604
rect 5194 1660 5258 1664
rect 5194 1604 5198 1660
rect 5198 1604 5254 1660
rect 5254 1604 5258 1660
rect 5194 1600 5258 1604
rect 5274 1660 5338 1664
rect 5274 1604 5278 1660
rect 5278 1604 5334 1660
rect 5334 1604 5338 1660
rect 5274 1600 5338 1604
rect 5354 1660 5418 1664
rect 5354 1604 5358 1660
rect 5358 1604 5414 1660
rect 5414 1604 5418 1660
rect 5354 1600 5418 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 10069 1660 10133 1664
rect 10069 1604 10073 1660
rect 10073 1604 10129 1660
rect 10129 1604 10133 1660
rect 10069 1600 10133 1604
rect 14544 1660 14608 1664
rect 14544 1604 14548 1660
rect 14548 1604 14604 1660
rect 14604 1604 14608 1660
rect 14544 1600 14608 1604
rect 14624 1660 14688 1664
rect 14624 1604 14628 1660
rect 14628 1604 14684 1660
rect 14684 1604 14688 1660
rect 14624 1600 14688 1604
rect 14704 1660 14768 1664
rect 14704 1604 14708 1660
rect 14708 1604 14764 1660
rect 14764 1604 14768 1660
rect 14704 1600 14768 1604
rect 14784 1660 14848 1664
rect 14784 1604 14788 1660
rect 14788 1604 14844 1660
rect 14844 1604 14848 1660
rect 14784 1600 14848 1604
rect 19259 1660 19323 1664
rect 19259 1604 19263 1660
rect 19263 1604 19319 1660
rect 19319 1604 19323 1660
rect 19259 1600 19323 1604
rect 19339 1660 19403 1664
rect 19339 1604 19343 1660
rect 19343 1604 19399 1660
rect 19399 1604 19403 1660
rect 19339 1600 19403 1604
rect 19419 1660 19483 1664
rect 19419 1604 19423 1660
rect 19423 1604 19479 1660
rect 19479 1604 19483 1660
rect 19419 1600 19483 1604
rect 19499 1660 19563 1664
rect 19499 1604 19503 1660
rect 19503 1604 19559 1660
rect 19559 1604 19563 1660
rect 19499 1600 19563 1604
rect 2757 1116 2821 1120
rect 2757 1060 2761 1116
rect 2761 1060 2817 1116
rect 2817 1060 2821 1116
rect 2757 1056 2821 1060
rect 2837 1116 2901 1120
rect 2837 1060 2841 1116
rect 2841 1060 2897 1116
rect 2897 1060 2901 1116
rect 2837 1056 2901 1060
rect 2917 1116 2981 1120
rect 2917 1060 2921 1116
rect 2921 1060 2977 1116
rect 2977 1060 2981 1116
rect 2917 1056 2981 1060
rect 2997 1116 3061 1120
rect 2997 1060 3001 1116
rect 3001 1060 3057 1116
rect 3057 1060 3061 1116
rect 2997 1056 3061 1060
rect 7472 1116 7536 1120
rect 7472 1060 7476 1116
rect 7476 1060 7532 1116
rect 7532 1060 7536 1116
rect 7472 1056 7536 1060
rect 7552 1116 7616 1120
rect 7552 1060 7556 1116
rect 7556 1060 7612 1116
rect 7612 1060 7616 1116
rect 7552 1056 7616 1060
rect 7632 1116 7696 1120
rect 7632 1060 7636 1116
rect 7636 1060 7692 1116
rect 7692 1060 7696 1116
rect 7632 1056 7696 1060
rect 7712 1116 7776 1120
rect 7712 1060 7716 1116
rect 7716 1060 7772 1116
rect 7772 1060 7776 1116
rect 7712 1056 7776 1060
rect 12187 1116 12251 1120
rect 12187 1060 12191 1116
rect 12191 1060 12247 1116
rect 12247 1060 12251 1116
rect 12187 1056 12251 1060
rect 12267 1116 12331 1120
rect 12267 1060 12271 1116
rect 12271 1060 12327 1116
rect 12327 1060 12331 1116
rect 12267 1056 12331 1060
rect 12347 1116 12411 1120
rect 12347 1060 12351 1116
rect 12351 1060 12407 1116
rect 12407 1060 12411 1116
rect 12347 1056 12411 1060
rect 12427 1116 12491 1120
rect 12427 1060 12431 1116
rect 12431 1060 12487 1116
rect 12487 1060 12491 1116
rect 12427 1056 12491 1060
rect 16902 1116 16966 1120
rect 16902 1060 16906 1116
rect 16906 1060 16962 1116
rect 16962 1060 16966 1116
rect 16902 1056 16966 1060
rect 16982 1116 17046 1120
rect 16982 1060 16986 1116
rect 16986 1060 17042 1116
rect 17042 1060 17046 1116
rect 16982 1056 17046 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 5114 572 5178 576
rect 5114 516 5118 572
rect 5118 516 5174 572
rect 5174 516 5178 572
rect 5114 512 5178 516
rect 5194 572 5258 576
rect 5194 516 5198 572
rect 5198 516 5254 572
rect 5254 516 5258 572
rect 5194 512 5258 516
rect 5274 572 5338 576
rect 5274 516 5278 572
rect 5278 516 5334 572
rect 5334 516 5338 572
rect 5274 512 5338 516
rect 5354 572 5418 576
rect 5354 516 5358 572
rect 5358 516 5414 572
rect 5414 516 5418 572
rect 5354 512 5418 516
rect 9829 572 9893 576
rect 9829 516 9833 572
rect 9833 516 9889 572
rect 9889 516 9893 572
rect 9829 512 9893 516
rect 9909 572 9973 576
rect 9909 516 9913 572
rect 9913 516 9969 572
rect 9969 516 9973 572
rect 9909 512 9973 516
rect 9989 572 10053 576
rect 9989 516 9993 572
rect 9993 516 10049 572
rect 10049 516 10053 572
rect 9989 512 10053 516
rect 10069 572 10133 576
rect 10069 516 10073 572
rect 10073 516 10129 572
rect 10129 516 10133 572
rect 10069 512 10133 516
rect 14544 572 14608 576
rect 14544 516 14548 572
rect 14548 516 14604 572
rect 14604 516 14608 572
rect 14544 512 14608 516
rect 14624 572 14688 576
rect 14624 516 14628 572
rect 14628 516 14684 572
rect 14684 516 14688 572
rect 14624 512 14688 516
rect 14704 572 14768 576
rect 14704 516 14708 572
rect 14708 516 14764 572
rect 14764 516 14768 572
rect 14704 512 14768 516
rect 14784 572 14848 576
rect 14784 516 14788 572
rect 14788 516 14844 572
rect 14844 516 14848 572
rect 14784 512 14848 516
rect 19259 572 19323 576
rect 19259 516 19263 572
rect 19263 516 19319 572
rect 19319 516 19323 572
rect 19259 512 19323 516
rect 19339 572 19403 576
rect 19339 516 19343 572
rect 19343 516 19399 572
rect 19399 516 19403 572
rect 19339 512 19403 516
rect 19419 572 19483 576
rect 19419 516 19423 572
rect 19423 516 19479 572
rect 19479 516 19483 572
rect 19419 512 19483 516
rect 19499 572 19563 576
rect 19499 516 19503 572
rect 19503 516 19559 572
rect 19559 516 19563 572
rect 19499 512 19563 516
<< metal4 >>
rect 2749 18528 3069 19088
rect 2749 18464 2757 18528
rect 2821 18464 2837 18528
rect 2901 18464 2917 18528
rect 2981 18464 2997 18528
rect 3061 18464 3069 18528
rect 2749 17440 3069 18464
rect 2749 17376 2757 17440
rect 2821 17376 2837 17440
rect 2901 17376 2917 17440
rect 2981 17376 2997 17440
rect 3061 17376 3069 17440
rect 2749 16352 3069 17376
rect 2749 16288 2757 16352
rect 2821 16288 2837 16352
rect 2901 16288 2917 16352
rect 2981 16288 2997 16352
rect 3061 16288 3069 16352
rect 2749 15264 3069 16288
rect 2749 15200 2757 15264
rect 2821 15200 2837 15264
rect 2901 15200 2917 15264
rect 2981 15200 2997 15264
rect 3061 15200 3069 15264
rect 2749 14176 3069 15200
rect 2749 14112 2757 14176
rect 2821 14112 2837 14176
rect 2901 14112 2917 14176
rect 2981 14112 2997 14176
rect 3061 14112 3069 14176
rect 2749 13088 3069 14112
rect 2749 13024 2757 13088
rect 2821 13024 2837 13088
rect 2901 13024 2917 13088
rect 2981 13024 2997 13088
rect 3061 13024 3069 13088
rect 2749 12000 3069 13024
rect 2749 11936 2757 12000
rect 2821 11936 2837 12000
rect 2901 11936 2917 12000
rect 2981 11936 2997 12000
rect 3061 11936 3069 12000
rect 2749 10912 3069 11936
rect 2749 10848 2757 10912
rect 2821 10848 2837 10912
rect 2901 10848 2917 10912
rect 2981 10848 2997 10912
rect 3061 10848 3069 10912
rect 2749 9824 3069 10848
rect 2749 9760 2757 9824
rect 2821 9760 2837 9824
rect 2901 9760 2917 9824
rect 2981 9760 2997 9824
rect 3061 9760 3069 9824
rect 2749 8736 3069 9760
rect 2749 8672 2757 8736
rect 2821 8672 2837 8736
rect 2901 8672 2917 8736
rect 2981 8672 2997 8736
rect 3061 8672 3069 8736
rect 2749 7648 3069 8672
rect 2749 7584 2757 7648
rect 2821 7584 2837 7648
rect 2901 7584 2917 7648
rect 2981 7584 2997 7648
rect 3061 7584 3069 7648
rect 2749 6560 3069 7584
rect 2749 6496 2757 6560
rect 2821 6496 2837 6560
rect 2901 6496 2917 6560
rect 2981 6496 2997 6560
rect 3061 6496 3069 6560
rect 2749 5472 3069 6496
rect 2749 5408 2757 5472
rect 2821 5408 2837 5472
rect 2901 5408 2917 5472
rect 2981 5408 2997 5472
rect 3061 5408 3069 5472
rect 2749 4384 3069 5408
rect 2749 4320 2757 4384
rect 2821 4320 2837 4384
rect 2901 4320 2917 4384
rect 2981 4320 2997 4384
rect 3061 4320 3069 4384
rect 2749 3296 3069 4320
rect 2749 3232 2757 3296
rect 2821 3232 2837 3296
rect 2901 3232 2917 3296
rect 2981 3232 2997 3296
rect 3061 3232 3069 3296
rect 2749 2208 3069 3232
rect 2749 2144 2757 2208
rect 2821 2144 2837 2208
rect 2901 2144 2917 2208
rect 2981 2144 2997 2208
rect 3061 2144 3069 2208
rect 2749 1120 3069 2144
rect 2749 1056 2757 1120
rect 2821 1056 2837 1120
rect 2901 1056 2917 1120
rect 2981 1056 2997 1120
rect 3061 1056 3069 1120
rect 2749 496 3069 1056
rect 5106 19072 5426 19088
rect 5106 19008 5114 19072
rect 5178 19008 5194 19072
rect 5258 19008 5274 19072
rect 5338 19008 5354 19072
rect 5418 19008 5426 19072
rect 5106 17984 5426 19008
rect 5106 17920 5114 17984
rect 5178 17920 5194 17984
rect 5258 17920 5274 17984
rect 5338 17920 5354 17984
rect 5418 17920 5426 17984
rect 5106 16896 5426 17920
rect 5106 16832 5114 16896
rect 5178 16832 5194 16896
rect 5258 16832 5274 16896
rect 5338 16832 5354 16896
rect 5418 16832 5426 16896
rect 5106 15808 5426 16832
rect 5106 15744 5114 15808
rect 5178 15744 5194 15808
rect 5258 15744 5274 15808
rect 5338 15744 5354 15808
rect 5418 15744 5426 15808
rect 5106 14720 5426 15744
rect 5106 14656 5114 14720
rect 5178 14656 5194 14720
rect 5258 14656 5274 14720
rect 5338 14656 5354 14720
rect 5418 14656 5426 14720
rect 5106 13632 5426 14656
rect 5106 13568 5114 13632
rect 5178 13568 5194 13632
rect 5258 13568 5274 13632
rect 5338 13568 5354 13632
rect 5418 13568 5426 13632
rect 5106 12544 5426 13568
rect 5106 12480 5114 12544
rect 5178 12480 5194 12544
rect 5258 12480 5274 12544
rect 5338 12480 5354 12544
rect 5418 12480 5426 12544
rect 5106 11456 5426 12480
rect 5106 11392 5114 11456
rect 5178 11392 5194 11456
rect 5258 11392 5274 11456
rect 5338 11392 5354 11456
rect 5418 11392 5426 11456
rect 5106 10368 5426 11392
rect 5106 10304 5114 10368
rect 5178 10304 5194 10368
rect 5258 10304 5274 10368
rect 5338 10304 5354 10368
rect 5418 10304 5426 10368
rect 5106 9280 5426 10304
rect 5106 9216 5114 9280
rect 5178 9216 5194 9280
rect 5258 9216 5274 9280
rect 5338 9216 5354 9280
rect 5418 9216 5426 9280
rect 5106 8192 5426 9216
rect 5106 8128 5114 8192
rect 5178 8128 5194 8192
rect 5258 8128 5274 8192
rect 5338 8128 5354 8192
rect 5418 8128 5426 8192
rect 5106 7104 5426 8128
rect 5106 7040 5114 7104
rect 5178 7040 5194 7104
rect 5258 7040 5274 7104
rect 5338 7040 5354 7104
rect 5418 7040 5426 7104
rect 5106 6016 5426 7040
rect 5106 5952 5114 6016
rect 5178 5952 5194 6016
rect 5258 5952 5274 6016
rect 5338 5952 5354 6016
rect 5418 5952 5426 6016
rect 5106 4928 5426 5952
rect 5106 4864 5114 4928
rect 5178 4864 5194 4928
rect 5258 4864 5274 4928
rect 5338 4864 5354 4928
rect 5418 4864 5426 4928
rect 5106 3840 5426 4864
rect 5106 3776 5114 3840
rect 5178 3776 5194 3840
rect 5258 3776 5274 3840
rect 5338 3776 5354 3840
rect 5418 3776 5426 3840
rect 5106 2752 5426 3776
rect 5106 2688 5114 2752
rect 5178 2688 5194 2752
rect 5258 2688 5274 2752
rect 5338 2688 5354 2752
rect 5418 2688 5426 2752
rect 5106 1664 5426 2688
rect 5106 1600 5114 1664
rect 5178 1600 5194 1664
rect 5258 1600 5274 1664
rect 5338 1600 5354 1664
rect 5418 1600 5426 1664
rect 5106 576 5426 1600
rect 5106 512 5114 576
rect 5178 512 5194 576
rect 5258 512 5274 576
rect 5338 512 5354 576
rect 5418 512 5426 576
rect 5106 496 5426 512
rect 7464 18528 7784 19088
rect 7464 18464 7472 18528
rect 7536 18464 7552 18528
rect 7616 18464 7632 18528
rect 7696 18464 7712 18528
rect 7776 18464 7784 18528
rect 7464 17440 7784 18464
rect 7464 17376 7472 17440
rect 7536 17376 7552 17440
rect 7616 17376 7632 17440
rect 7696 17376 7712 17440
rect 7776 17376 7784 17440
rect 7464 16352 7784 17376
rect 7464 16288 7472 16352
rect 7536 16288 7552 16352
rect 7616 16288 7632 16352
rect 7696 16288 7712 16352
rect 7776 16288 7784 16352
rect 7464 15264 7784 16288
rect 9821 19072 10141 19088
rect 9821 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10069 19072
rect 10133 19008 10141 19072
rect 9821 17984 10141 19008
rect 9821 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10069 17984
rect 10133 17920 10141 17984
rect 9821 16896 10141 17920
rect 9821 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10069 16896
rect 10133 16832 10141 16896
rect 9821 15808 10141 16832
rect 12179 18528 12499 19088
rect 12179 18464 12187 18528
rect 12251 18464 12267 18528
rect 12331 18464 12347 18528
rect 12411 18464 12427 18528
rect 12491 18464 12499 18528
rect 12179 17440 12499 18464
rect 12179 17376 12187 17440
rect 12251 17376 12267 17440
rect 12331 17376 12347 17440
rect 12411 17376 12427 17440
rect 12491 17376 12499 17440
rect 10363 16692 10429 16693
rect 10363 16628 10364 16692
rect 10428 16628 10429 16692
rect 10363 16627 10429 16628
rect 9821 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10069 15808
rect 10133 15744 10141 15808
rect 8707 15468 8773 15469
rect 8707 15404 8708 15468
rect 8772 15404 8773 15468
rect 8707 15403 8773 15404
rect 7464 15200 7472 15264
rect 7536 15200 7552 15264
rect 7616 15200 7632 15264
rect 7696 15200 7712 15264
rect 7776 15200 7784 15264
rect 7464 14176 7784 15200
rect 7464 14112 7472 14176
rect 7536 14112 7552 14176
rect 7616 14112 7632 14176
rect 7696 14112 7712 14176
rect 7776 14112 7784 14176
rect 7464 13088 7784 14112
rect 7464 13024 7472 13088
rect 7536 13024 7552 13088
rect 7616 13024 7632 13088
rect 7696 13024 7712 13088
rect 7776 13024 7784 13088
rect 7464 12000 7784 13024
rect 8710 12749 8770 15403
rect 9821 14720 10141 15744
rect 9821 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10069 14720
rect 10133 14656 10141 14720
rect 9821 13632 10141 14656
rect 9821 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10069 13632
rect 10133 13568 10141 13632
rect 8707 12748 8773 12749
rect 8707 12684 8708 12748
rect 8772 12684 8773 12748
rect 8707 12683 8773 12684
rect 7464 11936 7472 12000
rect 7536 11936 7552 12000
rect 7616 11936 7632 12000
rect 7696 11936 7712 12000
rect 7776 11936 7784 12000
rect 7464 10912 7784 11936
rect 7464 10848 7472 10912
rect 7536 10848 7552 10912
rect 7616 10848 7632 10912
rect 7696 10848 7712 10912
rect 7776 10848 7784 10912
rect 7464 9824 7784 10848
rect 7464 9760 7472 9824
rect 7536 9760 7552 9824
rect 7616 9760 7632 9824
rect 7696 9760 7712 9824
rect 7776 9760 7784 9824
rect 7464 8736 7784 9760
rect 7464 8672 7472 8736
rect 7536 8672 7552 8736
rect 7616 8672 7632 8736
rect 7696 8672 7712 8736
rect 7776 8672 7784 8736
rect 7464 7648 7784 8672
rect 7464 7584 7472 7648
rect 7536 7584 7552 7648
rect 7616 7584 7632 7648
rect 7696 7584 7712 7648
rect 7776 7584 7784 7648
rect 7464 6560 7784 7584
rect 7464 6496 7472 6560
rect 7536 6496 7552 6560
rect 7616 6496 7632 6560
rect 7696 6496 7712 6560
rect 7776 6496 7784 6560
rect 7464 5472 7784 6496
rect 7464 5408 7472 5472
rect 7536 5408 7552 5472
rect 7616 5408 7632 5472
rect 7696 5408 7712 5472
rect 7776 5408 7784 5472
rect 7464 4384 7784 5408
rect 7464 4320 7472 4384
rect 7536 4320 7552 4384
rect 7616 4320 7632 4384
rect 7696 4320 7712 4384
rect 7776 4320 7784 4384
rect 7464 3296 7784 4320
rect 7464 3232 7472 3296
rect 7536 3232 7552 3296
rect 7616 3232 7632 3296
rect 7696 3232 7712 3296
rect 7776 3232 7784 3296
rect 7464 2208 7784 3232
rect 7464 2144 7472 2208
rect 7536 2144 7552 2208
rect 7616 2144 7632 2208
rect 7696 2144 7712 2208
rect 7776 2144 7784 2208
rect 7464 1120 7784 2144
rect 7464 1056 7472 1120
rect 7536 1056 7552 1120
rect 7616 1056 7632 1120
rect 7696 1056 7712 1120
rect 7776 1056 7784 1120
rect 7464 496 7784 1056
rect 9821 12544 10141 13568
rect 9821 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10069 12544
rect 10133 12480 10141 12544
rect 9821 11456 10141 12480
rect 9821 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10069 11456
rect 10133 11392 10141 11456
rect 9821 10368 10141 11392
rect 9821 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10069 10368
rect 10133 10304 10141 10368
rect 9821 9280 10141 10304
rect 9821 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10069 9280
rect 10133 9216 10141 9280
rect 9821 8192 10141 9216
rect 9821 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10069 8192
rect 10133 8128 10141 8192
rect 9821 7104 10141 8128
rect 9821 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10069 7104
rect 10133 7040 10141 7104
rect 9821 6016 10141 7040
rect 10366 6901 10426 16627
rect 12179 16352 12499 17376
rect 12179 16288 12187 16352
rect 12251 16288 12267 16352
rect 12331 16288 12347 16352
rect 12411 16288 12427 16352
rect 12491 16288 12499 16352
rect 12179 15264 12499 16288
rect 12179 15200 12187 15264
rect 12251 15200 12267 15264
rect 12331 15200 12347 15264
rect 12411 15200 12427 15264
rect 12491 15200 12499 15264
rect 12179 14176 12499 15200
rect 12179 14112 12187 14176
rect 12251 14112 12267 14176
rect 12331 14112 12347 14176
rect 12411 14112 12427 14176
rect 12491 14112 12499 14176
rect 12179 13088 12499 14112
rect 12179 13024 12187 13088
rect 12251 13024 12267 13088
rect 12331 13024 12347 13088
rect 12411 13024 12427 13088
rect 12491 13024 12499 13088
rect 12179 12000 12499 13024
rect 12179 11936 12187 12000
rect 12251 11936 12267 12000
rect 12331 11936 12347 12000
rect 12411 11936 12427 12000
rect 12491 11936 12499 12000
rect 12179 10912 12499 11936
rect 12179 10848 12187 10912
rect 12251 10848 12267 10912
rect 12331 10848 12347 10912
rect 12411 10848 12427 10912
rect 12491 10848 12499 10912
rect 12179 9824 12499 10848
rect 12179 9760 12187 9824
rect 12251 9760 12267 9824
rect 12331 9760 12347 9824
rect 12411 9760 12427 9824
rect 12491 9760 12499 9824
rect 12179 8736 12499 9760
rect 12179 8672 12187 8736
rect 12251 8672 12267 8736
rect 12331 8672 12347 8736
rect 12411 8672 12427 8736
rect 12491 8672 12499 8736
rect 12179 7648 12499 8672
rect 12179 7584 12187 7648
rect 12251 7584 12267 7648
rect 12331 7584 12347 7648
rect 12411 7584 12427 7648
rect 12491 7584 12499 7648
rect 10363 6900 10429 6901
rect 10363 6836 10364 6900
rect 10428 6836 10429 6900
rect 10363 6835 10429 6836
rect 9821 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10069 6016
rect 10133 5952 10141 6016
rect 9821 4928 10141 5952
rect 9821 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10069 4928
rect 10133 4864 10141 4928
rect 9821 3840 10141 4864
rect 9821 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10069 3840
rect 10133 3776 10141 3840
rect 9821 2752 10141 3776
rect 9821 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10069 2752
rect 10133 2688 10141 2752
rect 9821 1664 10141 2688
rect 9821 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10069 1664
rect 10133 1600 10141 1664
rect 9821 576 10141 1600
rect 9821 512 9829 576
rect 9893 512 9909 576
rect 9973 512 9989 576
rect 10053 512 10069 576
rect 10133 512 10141 576
rect 9821 496 10141 512
rect 12179 6560 12499 7584
rect 12179 6496 12187 6560
rect 12251 6496 12267 6560
rect 12331 6496 12347 6560
rect 12411 6496 12427 6560
rect 12491 6496 12499 6560
rect 12179 5472 12499 6496
rect 12179 5408 12187 5472
rect 12251 5408 12267 5472
rect 12331 5408 12347 5472
rect 12411 5408 12427 5472
rect 12491 5408 12499 5472
rect 12179 4384 12499 5408
rect 12179 4320 12187 4384
rect 12251 4320 12267 4384
rect 12331 4320 12347 4384
rect 12411 4320 12427 4384
rect 12491 4320 12499 4384
rect 12179 3296 12499 4320
rect 12179 3232 12187 3296
rect 12251 3232 12267 3296
rect 12331 3232 12347 3296
rect 12411 3232 12427 3296
rect 12491 3232 12499 3296
rect 12179 2208 12499 3232
rect 12179 2144 12187 2208
rect 12251 2144 12267 2208
rect 12331 2144 12347 2208
rect 12411 2144 12427 2208
rect 12491 2144 12499 2208
rect 12179 1120 12499 2144
rect 12179 1056 12187 1120
rect 12251 1056 12267 1120
rect 12331 1056 12347 1120
rect 12411 1056 12427 1120
rect 12491 1056 12499 1120
rect 12179 496 12499 1056
rect 14536 19072 14856 19088
rect 14536 19008 14544 19072
rect 14608 19008 14624 19072
rect 14688 19008 14704 19072
rect 14768 19008 14784 19072
rect 14848 19008 14856 19072
rect 14536 17984 14856 19008
rect 14536 17920 14544 17984
rect 14608 17920 14624 17984
rect 14688 17920 14704 17984
rect 14768 17920 14784 17984
rect 14848 17920 14856 17984
rect 14536 16896 14856 17920
rect 14536 16832 14544 16896
rect 14608 16832 14624 16896
rect 14688 16832 14704 16896
rect 14768 16832 14784 16896
rect 14848 16832 14856 16896
rect 14536 15808 14856 16832
rect 14536 15744 14544 15808
rect 14608 15744 14624 15808
rect 14688 15744 14704 15808
rect 14768 15744 14784 15808
rect 14848 15744 14856 15808
rect 14536 14720 14856 15744
rect 14536 14656 14544 14720
rect 14608 14656 14624 14720
rect 14688 14656 14704 14720
rect 14768 14656 14784 14720
rect 14848 14656 14856 14720
rect 14536 13632 14856 14656
rect 14536 13568 14544 13632
rect 14608 13568 14624 13632
rect 14688 13568 14704 13632
rect 14768 13568 14784 13632
rect 14848 13568 14856 13632
rect 14536 12544 14856 13568
rect 14536 12480 14544 12544
rect 14608 12480 14624 12544
rect 14688 12480 14704 12544
rect 14768 12480 14784 12544
rect 14848 12480 14856 12544
rect 14536 11456 14856 12480
rect 14536 11392 14544 11456
rect 14608 11392 14624 11456
rect 14688 11392 14704 11456
rect 14768 11392 14784 11456
rect 14848 11392 14856 11456
rect 14536 10368 14856 11392
rect 14536 10304 14544 10368
rect 14608 10304 14624 10368
rect 14688 10304 14704 10368
rect 14768 10304 14784 10368
rect 14848 10304 14856 10368
rect 14536 9280 14856 10304
rect 14536 9216 14544 9280
rect 14608 9216 14624 9280
rect 14688 9216 14704 9280
rect 14768 9216 14784 9280
rect 14848 9216 14856 9280
rect 14536 8192 14856 9216
rect 14536 8128 14544 8192
rect 14608 8128 14624 8192
rect 14688 8128 14704 8192
rect 14768 8128 14784 8192
rect 14848 8128 14856 8192
rect 14536 7104 14856 8128
rect 14536 7040 14544 7104
rect 14608 7040 14624 7104
rect 14688 7040 14704 7104
rect 14768 7040 14784 7104
rect 14848 7040 14856 7104
rect 14536 6016 14856 7040
rect 14536 5952 14544 6016
rect 14608 5952 14624 6016
rect 14688 5952 14704 6016
rect 14768 5952 14784 6016
rect 14848 5952 14856 6016
rect 14536 4928 14856 5952
rect 14536 4864 14544 4928
rect 14608 4864 14624 4928
rect 14688 4864 14704 4928
rect 14768 4864 14784 4928
rect 14848 4864 14856 4928
rect 14536 3840 14856 4864
rect 14536 3776 14544 3840
rect 14608 3776 14624 3840
rect 14688 3776 14704 3840
rect 14768 3776 14784 3840
rect 14848 3776 14856 3840
rect 14536 2752 14856 3776
rect 14536 2688 14544 2752
rect 14608 2688 14624 2752
rect 14688 2688 14704 2752
rect 14768 2688 14784 2752
rect 14848 2688 14856 2752
rect 14536 1664 14856 2688
rect 14536 1600 14544 1664
rect 14608 1600 14624 1664
rect 14688 1600 14704 1664
rect 14768 1600 14784 1664
rect 14848 1600 14856 1664
rect 14536 576 14856 1600
rect 14536 512 14544 576
rect 14608 512 14624 576
rect 14688 512 14704 576
rect 14768 512 14784 576
rect 14848 512 14856 576
rect 14536 496 14856 512
rect 16894 18528 17214 19088
rect 16894 18464 16902 18528
rect 16966 18464 16982 18528
rect 17046 18464 17062 18528
rect 17126 18464 17142 18528
rect 17206 18464 17214 18528
rect 16894 17440 17214 18464
rect 16894 17376 16902 17440
rect 16966 17376 16982 17440
rect 17046 17376 17062 17440
rect 17126 17376 17142 17440
rect 17206 17376 17214 17440
rect 16894 16352 17214 17376
rect 16894 16288 16902 16352
rect 16966 16288 16982 16352
rect 17046 16288 17062 16352
rect 17126 16288 17142 16352
rect 17206 16288 17214 16352
rect 16894 15264 17214 16288
rect 19251 19072 19571 19088
rect 19251 19008 19259 19072
rect 19323 19008 19339 19072
rect 19403 19008 19419 19072
rect 19483 19008 19499 19072
rect 19563 19008 19571 19072
rect 19251 17984 19571 19008
rect 19251 17920 19259 17984
rect 19323 17920 19339 17984
rect 19403 17920 19419 17984
rect 19483 17920 19499 17984
rect 19563 17920 19571 17984
rect 19251 16896 19571 17920
rect 19251 16832 19259 16896
rect 19323 16832 19339 16896
rect 19403 16832 19419 16896
rect 19483 16832 19499 16896
rect 19563 16832 19571 16896
rect 17907 16012 17973 16013
rect 17907 15948 17908 16012
rect 17972 15948 17973 16012
rect 17907 15947 17973 15948
rect 16894 15200 16902 15264
rect 16966 15200 16982 15264
rect 17046 15200 17062 15264
rect 17126 15200 17142 15264
rect 17206 15200 17214 15264
rect 16894 14176 17214 15200
rect 16894 14112 16902 14176
rect 16966 14112 16982 14176
rect 17046 14112 17062 14176
rect 17126 14112 17142 14176
rect 17206 14112 17214 14176
rect 16894 13088 17214 14112
rect 16894 13024 16902 13088
rect 16966 13024 16982 13088
rect 17046 13024 17062 13088
rect 17126 13024 17142 13088
rect 17206 13024 17214 13088
rect 16894 12000 17214 13024
rect 16894 11936 16902 12000
rect 16966 11936 16982 12000
rect 17046 11936 17062 12000
rect 17126 11936 17142 12000
rect 17206 11936 17214 12000
rect 16894 10912 17214 11936
rect 17910 11797 17970 15947
rect 19251 15808 19571 16832
rect 19251 15744 19259 15808
rect 19323 15744 19339 15808
rect 19403 15744 19419 15808
rect 19483 15744 19499 15808
rect 19563 15744 19571 15808
rect 19251 14720 19571 15744
rect 19251 14656 19259 14720
rect 19323 14656 19339 14720
rect 19403 14656 19419 14720
rect 19483 14656 19499 14720
rect 19563 14656 19571 14720
rect 19251 13632 19571 14656
rect 19251 13568 19259 13632
rect 19323 13568 19339 13632
rect 19403 13568 19419 13632
rect 19483 13568 19499 13632
rect 19563 13568 19571 13632
rect 19251 12544 19571 13568
rect 19251 12480 19259 12544
rect 19323 12480 19339 12544
rect 19403 12480 19419 12544
rect 19483 12480 19499 12544
rect 19563 12480 19571 12544
rect 17907 11796 17973 11797
rect 17907 11732 17908 11796
rect 17972 11732 17973 11796
rect 17907 11731 17973 11732
rect 16894 10848 16902 10912
rect 16966 10848 16982 10912
rect 17046 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17214 10912
rect 16894 9824 17214 10848
rect 16894 9760 16902 9824
rect 16966 9760 16982 9824
rect 17046 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17214 9824
rect 16894 8736 17214 9760
rect 16894 8672 16902 8736
rect 16966 8672 16982 8736
rect 17046 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17214 8736
rect 16894 7648 17214 8672
rect 16894 7584 16902 7648
rect 16966 7584 16982 7648
rect 17046 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17214 7648
rect 16894 6560 17214 7584
rect 16894 6496 16902 6560
rect 16966 6496 16982 6560
rect 17046 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17214 6560
rect 16894 5472 17214 6496
rect 16894 5408 16902 5472
rect 16966 5408 16982 5472
rect 17046 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17214 5472
rect 16894 4384 17214 5408
rect 16894 4320 16902 4384
rect 16966 4320 16982 4384
rect 17046 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17214 4384
rect 16894 3296 17214 4320
rect 16894 3232 16902 3296
rect 16966 3232 16982 3296
rect 17046 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17214 3296
rect 16894 2208 17214 3232
rect 16894 2144 16902 2208
rect 16966 2144 16982 2208
rect 17046 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17214 2208
rect 16894 1120 17214 2144
rect 16894 1056 16902 1120
rect 16966 1056 16982 1120
rect 17046 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17214 1120
rect 16894 496 17214 1056
rect 19251 11456 19571 12480
rect 19251 11392 19259 11456
rect 19323 11392 19339 11456
rect 19403 11392 19419 11456
rect 19483 11392 19499 11456
rect 19563 11392 19571 11456
rect 19251 10368 19571 11392
rect 19251 10304 19259 10368
rect 19323 10304 19339 10368
rect 19403 10304 19419 10368
rect 19483 10304 19499 10368
rect 19563 10304 19571 10368
rect 19251 9280 19571 10304
rect 19251 9216 19259 9280
rect 19323 9216 19339 9280
rect 19403 9216 19419 9280
rect 19483 9216 19499 9280
rect 19563 9216 19571 9280
rect 19251 8192 19571 9216
rect 19251 8128 19259 8192
rect 19323 8128 19339 8192
rect 19403 8128 19419 8192
rect 19483 8128 19499 8192
rect 19563 8128 19571 8192
rect 19251 7104 19571 8128
rect 19251 7040 19259 7104
rect 19323 7040 19339 7104
rect 19403 7040 19419 7104
rect 19483 7040 19499 7104
rect 19563 7040 19571 7104
rect 19251 6016 19571 7040
rect 19251 5952 19259 6016
rect 19323 5952 19339 6016
rect 19403 5952 19419 6016
rect 19483 5952 19499 6016
rect 19563 5952 19571 6016
rect 19251 4928 19571 5952
rect 19251 4864 19259 4928
rect 19323 4864 19339 4928
rect 19403 4864 19419 4928
rect 19483 4864 19499 4928
rect 19563 4864 19571 4928
rect 19251 3840 19571 4864
rect 19251 3776 19259 3840
rect 19323 3776 19339 3840
rect 19403 3776 19419 3840
rect 19483 3776 19499 3840
rect 19563 3776 19571 3840
rect 19251 2752 19571 3776
rect 19251 2688 19259 2752
rect 19323 2688 19339 2752
rect 19403 2688 19419 2752
rect 19483 2688 19499 2752
rect 19563 2688 19571 2752
rect 19251 1664 19571 2688
rect 19251 1600 19259 1664
rect 19323 1600 19339 1664
rect 19403 1600 19419 1664
rect 19483 1600 19499 1664
rect 19563 1600 19571 1664
rect 19251 576 19571 1600
rect 19251 512 19259 576
rect 19323 512 19339 576
rect 19403 512 19419 576
rect 19483 512 19499 576
rect 19563 512 19571 576
rect 19251 496 19571 512
use sky130_fd_sc_hd__inv_2  _212_
timestamp -3600
transform -1 0 4140 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _213_
timestamp -3600
transform -1 0 8832 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _214_
timestamp -3600
transform -1 0 8188 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _215_
timestamp -3600
transform 1 0 3956 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _216_
timestamp -3600
transform 1 0 6348 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _217_
timestamp -3600
transform 1 0 7452 0 -1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _218_
timestamp -3600
transform 1 0 4232 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp -3600
transform -1 0 6716 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp -3600
transform 1 0 11316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _221_
timestamp -3600
transform 1 0 4140 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _222_
timestamp -3600
transform 1 0 4876 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp -3600
transform 1 0 10672 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _224_
timestamp -3600
transform 1 0 4876 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _225_
timestamp -3600
transform 1 0 5612 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _226_
timestamp -3600
transform 1 0 5796 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor4b_1  _227_
timestamp -3600
transform -1 0 5704 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _228_
timestamp -3600
transform 1 0 10948 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _229_
timestamp -3600
transform 1 0 11408 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _230_
timestamp -3600
transform -1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _231_
timestamp -3600
transform -1 0 3956 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _232_
timestamp -3600
transform 1 0 3404 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _233_
timestamp -3600
transform 1 0 2024 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _234_
timestamp -3600
transform -1 0 2024 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _235_
timestamp -3600
transform -1 0 2944 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _236_
timestamp -3600
transform 1 0 2300 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _237_
timestamp -3600
transform -1 0 2392 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _238_
timestamp -3600
transform 1 0 1656 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _239_
timestamp -3600
transform -1 0 1748 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _240_
timestamp -3600
transform -1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _241_
timestamp -3600
transform 1 0 1748 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _242_
timestamp -3600
transform 1 0 2484 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _243_
timestamp -3600
transform 1 0 2484 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _244_
timestamp -3600
transform -1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _245_
timestamp -3600
transform 1 0 4048 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _246_
timestamp -3600
transform 1 0 3588 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _247_
timestamp -3600
transform -1 0 4600 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp -3600
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _249_
timestamp -3600
transform 1 0 4784 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp -3600
transform 1 0 4692 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _251_
timestamp -3600
transform 1 0 4876 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp -3600
transform -1 0 5612 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _253_
timestamp -3600
transform 1 0 5796 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _254_
timestamp -3600
transform 1 0 4692 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _255_
timestamp -3600
transform 1 0 5060 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp -3600
transform 1 0 6992 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _257_
timestamp -3600
transform -1 0 5888 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp -3600
transform -1 0 6164 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _259_
timestamp -3600
transform 1 0 4968 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _260_
timestamp -3600
transform -1 0 6716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _261_
timestamp -3600
transform -1 0 4968 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _262_
timestamp -3600
transform 1 0 4416 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _263_
timestamp -3600
transform 1 0 3680 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp -3600
transform 1 0 3956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _265_
timestamp -3600
transform 1 0 2300 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _266_
timestamp -3600
transform -1 0 3220 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _267_
timestamp -3600
transform -1 0 2760 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _268_
timestamp -3600
transform 1 0 1840 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _269_
timestamp -3600
transform -1 0 2852 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _270_
timestamp -3600
transform -1 0 3220 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _271_
timestamp -3600
transform -1 0 2944 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _272_
timestamp -3600
transform -1 0 3036 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _273_
timestamp -3600
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _274_
timestamp -3600
transform 1 0 7544 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _275_
timestamp -3600
transform 1 0 10212 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp -3600
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _277_
timestamp -3600
transform -1 0 10212 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _278_
timestamp -3600
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  _279_
timestamp -3600
transform -1 0 14352 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _280_
timestamp -3600
transform 1 0 10948 0 -1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _281_
timestamp -3600
transform 1 0 12880 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _282_
timestamp -3600
transform 1 0 16928 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _283_
timestamp -3600
transform 1 0 16100 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _284_
timestamp -3600
transform 1 0 13984 0 -1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _285_
timestamp -3600
transform 1 0 18308 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _286_
timestamp -3600
transform 1 0 13984 0 -1 14688
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  _287_
timestamp -3600
transform 1 0 17480 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _288_
timestamp -3600
transform -1 0 17020 0 1 13600
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _289_
timestamp -3600
transform -1 0 16744 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _290_
timestamp -3600
transform 1 0 16744 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _291_
timestamp -3600
transform 1 0 11224 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _292_
timestamp -3600
transform 1 0 12420 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _293_
timestamp -3600
transform 1 0 16744 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_4  _294_
timestamp -3600
transform 1 0 14352 0 1 12512
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _295_
timestamp -3600
transform -1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _296_
timestamp -3600
transform -1 0 16008 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _297_
timestamp -3600
transform -1 0 16008 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _298_
timestamp -3600
transform 1 0 11224 0 -1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__a211o_1  _299_
timestamp -3600
transform 1 0 15548 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _300_
timestamp -3600
transform 1 0 17388 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _301_
timestamp -3600
transform -1 0 16744 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _302_
timestamp -3600
transform 1 0 16100 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _303_
timestamp -3600
transform 1 0 15640 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _304_
timestamp -3600
transform 1 0 14904 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _305_
timestamp -3600
transform 1 0 8464 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _306_
timestamp -3600
transform -1 0 11684 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _307_
timestamp -3600
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _308_
timestamp -3600
transform -1 0 8740 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _309_
timestamp -3600
transform 1 0 9200 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _310_
timestamp -3600
transform 1 0 13524 0 1 11424
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _311_
timestamp -3600
transform 1 0 14352 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _312_
timestamp -3600
transform 1 0 16008 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _313_
timestamp -3600
transform 1 0 16100 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _314_
timestamp -3600
transform 1 0 15732 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _315_
timestamp -3600
transform 1 0 16468 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _316_
timestamp -3600
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _317_
timestamp -3600
transform 1 0 15456 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _318_
timestamp -3600
transform 1 0 16100 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _319_
timestamp -3600
transform -1 0 17204 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _320_
timestamp -3600
transform -1 0 15916 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _321_
timestamp -3600
transform 1 0 14444 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _322_
timestamp -3600
transform 1 0 14996 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _323_
timestamp -3600
transform -1 0 14628 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _324_
timestamp -3600
transform 1 0 14996 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _325_
timestamp -3600
transform 1 0 8832 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _326_
timestamp -3600
transform 1 0 8464 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _327_
timestamp -3600
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _328_
timestamp -3600
transform 1 0 10764 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _329_
timestamp -3600
transform 1 0 15180 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _330_
timestamp -3600
transform 1 0 13984 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _331_
timestamp -3600
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _332_
timestamp -3600
transform 1 0 14076 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _333_
timestamp -3600
transform 1 0 16100 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _334_
timestamp -3600
transform 1 0 14628 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp -3600
transform -1 0 14076 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _336_
timestamp -3600
transform 1 0 14260 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _337_
timestamp -3600
transform 1 0 13708 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _338_
timestamp -3600
transform -1 0 14812 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _339_
timestamp -3600
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _340_
timestamp -3600
transform 1 0 13708 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _341_
timestamp -3600
transform 1 0 12972 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp -3600
transform 1 0 8464 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _343_
timestamp -3600
transform -1 0 7728 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _344_
timestamp -3600
transform -1 0 13800 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _345_
timestamp -3600
transform -1 0 14168 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _346_
timestamp -3600
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _347_
timestamp -3600
transform 1 0 12972 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _348_
timestamp -3600
transform 1 0 12236 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _349_
timestamp -3600
transform -1 0 13984 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _350_
timestamp -3600
transform 1 0 11592 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _351_
timestamp -3600
transform -1 0 18216 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _352_
timestamp -3600
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _353_
timestamp -3600
transform -1 0 13432 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _354_
timestamp -3600
transform 1 0 12788 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _355_
timestamp -3600
transform -1 0 12512 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _356_
timestamp -3600
transform 1 0 10028 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _357_
timestamp -3600
transform -1 0 10672 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _358_
timestamp -3600
transform 1 0 9292 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _359_
timestamp -3600
transform 1 0 8832 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _360_
timestamp -3600
transform -1 0 9752 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _361_
timestamp -3600
transform 1 0 12236 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _362_
timestamp -3600
transform -1 0 13800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp -3600
transform -1 0 11776 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _364_
timestamp -3600
transform 1 0 13708 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _365_
timestamp -3600
transform -1 0 13432 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _366_
timestamp -3600
transform 1 0 11776 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp -3600
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _368_
timestamp -3600
transform -1 0 10304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _369_
timestamp -3600
transform -1 0 10120 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp -3600
transform -1 0 13064 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _371_
timestamp -3600
transform -1 0 13156 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _372_
timestamp -3600
transform -1 0 11132 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _373_
timestamp -3600
transform -1 0 11316 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _374_
timestamp -3600
transform -1 0 7176 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp -3600
transform -1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _376_
timestamp -3600
transform -1 0 10672 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _377_
timestamp -3600
transform -1 0 10856 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _378_
timestamp -3600
transform -1 0 10396 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _379_
timestamp -3600
transform -1 0 16836 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _380_
timestamp -3600
transform 1 0 11408 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _381_
timestamp -3600
transform -1 0 11868 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _382_
timestamp -3600
transform 1 0 12052 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _383_
timestamp -3600
transform 1 0 11776 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _384_
timestamp -3600
transform 1 0 11316 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp -3600
transform -1 0 13156 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _386_
timestamp -3600
transform -1 0 14076 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _387_
timestamp -3600
transform 1 0 11960 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _388_
timestamp -3600
transform -1 0 12972 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp -3600
transform -1 0 12880 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _390_
timestamp -3600
transform 1 0 11684 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _391_
timestamp -3600
transform 1 0 11592 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _392_
timestamp -3600
transform 1 0 11684 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp -3600
transform -1 0 11408 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _394_
timestamp -3600
transform -1 0 11500 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _395_
timestamp -3600
transform -1 0 10120 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _396_
timestamp -3600
transform 1 0 9936 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _397_
timestamp -3600
transform 1 0 9476 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _398_
timestamp -3600
transform 1 0 8464 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _399_
timestamp -3600
transform -1 0 10856 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _400_
timestamp -3600
transform -1 0 10856 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _401_
timestamp -3600
transform -1 0 10948 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _402_
timestamp -3600
transform -1 0 8464 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _403_
timestamp -3600
transform -1 0 10028 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _404_
timestamp -3600
transform -1 0 10488 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp -3600
transform 1 0 9016 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _406_
timestamp -3600
transform 1 0 8280 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _407_
timestamp -3600
transform 1 0 6716 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _408_
timestamp -3600
transform 1 0 7176 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _409_
timestamp -3600
transform -1 0 9476 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _410_
timestamp -3600
transform 1 0 9108 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _411_
timestamp -3600
transform 1 0 7268 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _412_
timestamp -3600
transform -1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _413_
timestamp -3600
transform 1 0 9752 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _414_
timestamp -3600
transform 1 0 9384 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _415_
timestamp -3600
transform 1 0 7912 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _416_
timestamp -3600
transform 1 0 8372 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _417_
timestamp -3600
transform 1 0 8648 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _418_
timestamp -3600
transform 1 0 9108 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _419_
timestamp -3600
transform -1 0 6808 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _420_
timestamp -3600
transform -1 0 6808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _421_
timestamp -3600
transform -1 0 9108 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _422_
timestamp -3600
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _423_
timestamp -3600
transform 1 0 3036 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _424_
timestamp -3600
transform 1 0 1564 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _425_
timestamp -3600
transform 1 0 828 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _426_
timestamp -3600
transform -1 0 3864 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _427_
timestamp -3600
transform -1 0 4784 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _428_
timestamp -3600
transform -1 0 7268 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _429_
timestamp -3600
transform -1 0 7268 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _430_
timestamp -3600
transform 1 0 6256 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _431_
timestamp -3600
transform 1 0 3496 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _432_
timestamp -3600
transform 1 0 1656 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _433_
timestamp -3600
transform 1 0 1196 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _434_
timestamp -3600
transform 1 0 1012 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _435_
timestamp -3600
transform -1 0 8280 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _436_
timestamp -3600
transform -1 0 9936 0 1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _437_
timestamp -3600
transform -1 0 8004 0 1 9248
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _438_
timestamp -3600
transform -1 0 9936 0 1 8160
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _439_
timestamp -3600
transform 1 0 9292 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _440_
timestamp -3600
transform 1 0 11132 0 1 4896
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _441_
timestamp -3600
transform 1 0 10948 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _442_
timestamp -3600
transform 1 0 16744 0 -1 5984
box -38 -48 1602 592
use sky130_fd_sc_hd__conb_1  _443__15
timestamp -3600
transform 1 0 14904 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _443_
timestamp -3600
transform 1 0 14168 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_2  _444_
timestamp -3600
transform 1 0 11868 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _445_
timestamp -3600
transform 1 0 13524 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _446_
timestamp -3600
transform 1 0 12420 0 -1 14688
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _447_
timestamp -3600
transform 1 0 12052 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _448_
timestamp -3600
transform 1 0 9292 0 -1 13600
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _449_
timestamp -3600
transform 1 0 7728 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _450_
timestamp -3600
transform 1 0 10948 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _451_
timestamp -3600
transform 1 0 8372 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _452_
timestamp -3600
transform -1 0 8188 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _453_
timestamp -3600
transform 1 0 9844 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _454_
timestamp -3600
transform 1 0 6256 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _455_
timestamp -3600
transform 1 0 9108 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _456_
timestamp -3600
transform -1 0 8280 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _457_
timestamp -3600
transform 1 0 9200 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _458_
timestamp -3600
transform -1 0 5888 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _459_
timestamp -3600
transform -1 0 9844 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -3600
transform -1 0 10672 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -3600
transform -1 0 6992 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -3600
transform -1 0 8740 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -3600
transform 1 0 10396 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -3600
transform 1 0 11500 0 1 12512
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp -3600
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp -3600
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp -3600
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp -3600
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp -3600
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp -3600
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp -3600
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp -3600
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp -3600
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp -3600
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp -3600
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp -3600
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp -3600
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp -3600
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp -3600
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp -3600
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp -3600
transform 1 0 14628 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp -3600
transform 1 0 15732 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp -3600
transform 1 0 16100 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp -3600
transform 1 0 17204 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp -3600
transform 1 0 18308 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197
timestamp -3600
transform 1 0 18676 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_201
timestamp -3600
transform 1 0 19044 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp -3600
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp -3600
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp -3600
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp -3600
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp -3600
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp -3600
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp -3600
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp -3600
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp -3600
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp -3600
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp -3600
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp -3600
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp -3600
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp -3600
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp -3600
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp -3600
transform 1 0 14260 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp -3600
transform 1 0 15364 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp -3600
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp -3600
transform 1 0 16100 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp -3600
transform 1 0 17204 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_193
timestamp -3600
transform 1 0 18308 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_201
timestamp -3600
transform 1 0 19044 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp -3600
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp -3600
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp -3600
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp -3600
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp -3600
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp -3600
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp -3600
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp -3600
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp -3600
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp -3600
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp -3600
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp -3600
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp -3600
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp -3600
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp -3600
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp -3600
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp -3600
transform 1 0 14628 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp -3600
transform 1 0 15732 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp -3600
transform 1 0 16836 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp -3600
transform 1 0 17940 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp -3600
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp -3600
transform 1 0 18676 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp -3600
transform 1 0 19044 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp -3600
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp -3600
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp -3600
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp -3600
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp -3600
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp -3600
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp -3600
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp -3600
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp -3600
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp -3600
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp -3600
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp -3600
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp -3600
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp -3600
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp -3600
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp -3600
transform 1 0 14260 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp -3600
transform 1 0 15364 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp -3600
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp -3600
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp -3600
transform 1 0 17204 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_193
timestamp -3600
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp -3600
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp -3600
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp -3600
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp -3600
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp -3600
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp -3600
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp -3600
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp -3600
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp -3600
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp -3600
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp -3600
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp -3600
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp -3600
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp -3600
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp -3600
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp -3600
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp -3600
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp -3600
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp -3600
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp -3600
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp -3600
transform 1 0 17940 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp -3600
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_197
timestamp -3600
transform 1 0 18676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_201
timestamp -3600
transform 1 0 19044 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp -3600
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp -3600
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp -3600
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp -3600
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp -3600
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp -3600
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp -3600
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp -3600
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp -3600
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp -3600
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp -3600
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp -3600
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp -3600
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp -3600
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp -3600
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp -3600
transform 1 0 14260 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp -3600
transform 1 0 15364 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp -3600
transform 1 0 15916 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp -3600
transform 1 0 16100 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp -3600
transform 1 0 17204 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp -3600
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_201
timestamp -3600
transform 1 0 19044 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp -3600
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp -3600
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp -3600
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp -3600
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp -3600
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp -3600
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp -3600
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp -3600
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp -3600
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp -3600
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp -3600
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp -3600
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp -3600
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp -3600
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp -3600
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp -3600
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp -3600
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp -3600
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp -3600
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp -3600
transform 1 0 17940 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp -3600
transform 1 0 18492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp -3600
transform 1 0 18676 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp -3600
transform 1 0 19044 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp -3600
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp -3600
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp -3600
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp -3600
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp -3600
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp -3600
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp -3600
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp -3600
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp -3600
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp -3600
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp -3600
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp -3600
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp -3600
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp -3600
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp -3600
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp -3600
transform 1 0 14260 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp -3600
transform 1 0 15364 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp -3600
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp -3600
transform 1 0 16100 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp -3600
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp -3600
transform 1 0 18308 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_201
timestamp -3600
transform 1 0 19044 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp -3600
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp -3600
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp -3600
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp -3600
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp -3600
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp -3600
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp -3600
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp -3600
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp -3600
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp -3600
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp -3600
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_109
timestamp -3600
transform 1 0 10580 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_132
timestamp -3600
transform 1 0 12696 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp -3600
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp -3600
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp -3600
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp -3600
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp -3600
transform 1 0 17940 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp -3600
transform 1 0 18492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_197
timestamp -3600
transform 1 0 18676 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_201
timestamp -3600
transform 1 0 19044 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp -3600
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp -3600
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp -3600
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp -3600
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp -3600
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp -3600
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp -3600
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp -3600
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp -3600
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_93
timestamp -3600
transform 1 0 9108 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_130
timestamp -3600
transform 1 0 12512 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_142
timestamp -3600
transform 1 0 13616 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_154
timestamp -3600
transform 1 0 14720 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp -3600
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp -3600
transform 1 0 16100 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_175
timestamp -3600
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_193
timestamp -3600
transform 1 0 18308 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_201
timestamp -3600
transform 1 0 19044 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp -3600
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp -3600
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp -3600
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp -3600
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp -3600
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp -3600
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp -3600
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp -3600
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp -3600
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_110
timestamp -3600
transform 1 0 10672 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_122
timestamp -3600
transform 1 0 11776 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp -3600
transform 1 0 12880 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp -3600
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp -3600
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp -3600
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp -3600
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp -3600
transform 1 0 17940 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp -3600
transform 1 0 18492 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp -3600
transform 1 0 18676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp -3600
transform 1 0 19044 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp -3600
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp -3600
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp -3600
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp -3600
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp -3600
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp -3600
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp -3600
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp -3600
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_81
timestamp -3600
transform 1 0 8004 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_85
timestamp -3600
transform 1 0 8372 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_99
timestamp -3600
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp -3600
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_117
timestamp -3600
transform 1 0 11316 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_125
timestamp -3600
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_136
timestamp -3600
transform 1 0 13064 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_140
timestamp -3600
transform 1 0 13432 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_144
timestamp -3600
transform 1 0 13800 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_148
timestamp -3600
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_153
timestamp -3600
transform 1 0 14628 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_165
timestamp -3600
transform 1 0 15732 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_173
timestamp -3600
transform 1 0 16468 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_185
timestamp -3600
transform 1 0 17572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_197
timestamp -3600
transform 1 0 18676 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_201
timestamp -3600
transform 1 0 19044 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp -3600
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp -3600
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp -3600
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp -3600
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp -3600
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp -3600
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_89
timestamp -3600
transform 1 0 8740 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_115
timestamp -3600
transform 1 0 11132 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp -3600
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_161
timestamp -3600
transform 1 0 15364 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_167
timestamp -3600
transform 1 0 15916 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_179
timestamp -3600
transform 1 0 17020 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_191
timestamp -3600
transform 1 0 18124 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp -3600
transform 1 0 18492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp -3600
transform 1 0 18676 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp -3600
transform 1 0 19044 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp -3600
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp -3600
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp -3600
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp -3600
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp -3600
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp -3600
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp -3600
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp -3600
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_81
timestamp -3600
transform 1 0 8004 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp -3600
transform 1 0 8372 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_95
timestamp -3600
transform 1 0 9292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp -3600
transform 1 0 10396 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp -3600
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp -3600
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp -3600
transform 1 0 12052 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_133
timestamp -3600
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_141
timestamp -3600
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_149
timestamp -3600
transform 1 0 14260 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_155
timestamp -3600
transform 1 0 14812 0 -1 8160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_180
timestamp -3600
transform 1 0 17112 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_192
timestamp -3600
transform 1 0 18216 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_200
timestamp -3600
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp -3600
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp -3600
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp -3600
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp -3600
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp -3600
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp -3600
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp -3600
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp -3600
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp -3600
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_102
timestamp -3600
transform 1 0 9936 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_106
timestamp -3600
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_133
timestamp -3600
transform 1 0 12788 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp -3600
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_155
timestamp -3600
transform 1 0 14812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_170
timestamp -3600
transform 1 0 16192 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp -3600
transform 1 0 18676 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp -3600
transform 1 0 19044 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp -3600
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp -3600
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp -3600
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp -3600
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp -3600
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp -3600
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp -3600
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp -3600
transform 1 0 6900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_73
timestamp -3600
transform 1 0 7268 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_78
timestamp -3600
transform 1 0 7728 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_94
timestamp -3600
transform 1 0 9200 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp -3600
transform 1 0 10580 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp -3600
transform 1 0 10948 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp -3600
transform 1 0 11500 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_130
timestamp -3600
transform 1 0 12512 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_142
timestamp -3600
transform 1 0 13616 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_154
timestamp -3600
transform 1 0 14720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_162
timestamp -3600
transform 1 0 15456 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_176
timestamp -3600
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_192
timestamp -3600
transform 1 0 18216 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_200
timestamp -3600
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp -3600
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp -3600
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp -3600
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp -3600
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp -3600
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_53
timestamp -3600
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_61
timestamp -3600
transform 1 0 6164 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp -3600
transform 1 0 8004 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_85
timestamp -3600
transform 1 0 8372 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_95
timestamp -3600
transform 1 0 9292 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_110
timestamp -3600
transform 1 0 10672 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_124
timestamp -3600
transform 1 0 11960 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp -3600
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_149
timestamp -3600
transform 1 0 14260 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_161
timestamp -3600
transform 1 0 15364 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_173
timestamp -3600
transform 1 0 16468 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_185
timestamp -3600
transform 1 0 17572 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp -3600
transform 1 0 18308 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp -3600
transform 1 0 18676 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_201
timestamp -3600
transform 1 0 19044 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp -3600
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp -3600
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp -3600
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp -3600
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp -3600
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp -3600
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp -3600
transform 1 0 5796 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_72
timestamp -3600
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_77
timestamp -3600
transform 1 0 7636 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_89
timestamp -3600
transform 1 0 8740 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_97
timestamp -3600
transform 1 0 9476 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp -3600
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_155
timestamp -3600
transform 1 0 14812 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp -3600
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_173
timestamp -3600
transform 1 0 16468 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_181
timestamp -3600
transform 1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_192
timestamp -3600
transform 1 0 18216 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_200
timestamp -3600
transform 1 0 18952 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp -3600
transform 1 0 828 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp -3600
transform 1 0 1564 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp -3600
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp -3600
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp -3600
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_65
timestamp -3600
transform 1 0 6532 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_73
timestamp -3600
transform 1 0 7268 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp -3600
transform 1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp -3600
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_101
timestamp -3600
transform 1 0 9844 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_113
timestamp -3600
transform 1 0 10948 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_123
timestamp -3600
transform 1 0 11868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp -3600
transform 1 0 12972 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp -3600
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_160
timestamp -3600
transform 1 0 15272 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_164
timestamp -3600
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_177
timestamp -3600
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_182
timestamp -3600
transform 1 0 17296 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp -3600
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp -3600
transform 1 0 18676 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp -3600
transform 1 0 19044 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_3
timestamp -3600
transform 1 0 828 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_11
timestamp -3600
transform 1 0 1564 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_29
timestamp -3600
transform 1 0 3220 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_33
timestamp -3600
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_41
timestamp -3600
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp -3600
transform 1 0 4968 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp -3600
transform 1 0 5796 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_63
timestamp -3600
transform 1 0 6348 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_67
timestamp -3600
transform 1 0 6716 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_79
timestamp -3600
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_95
timestamp -3600
transform 1 0 9292 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_108
timestamp -3600
transform 1 0 10488 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp -3600
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_138
timestamp -3600
transform 1 0 13248 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_149
timestamp -3600
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_159
timestamp -3600
transform 1 0 15180 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp -3600
transform 1 0 17204 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_193
timestamp -3600
transform 1 0 18308 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp -3600
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp -3600
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_15
timestamp -3600
transform 1 0 1932 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp -3600
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp -3600
transform 1 0 3220 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_61
timestamp -3600
transform 1 0 6164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_78
timestamp -3600
transform 1 0 7728 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp -3600
transform 1 0 8372 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp -3600
transform 1 0 8740 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_113
timestamp -3600
transform 1 0 10948 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_125
timestamp -3600
transform 1 0 12052 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp -3600
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_154
timestamp -3600
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_158
timestamp -3600
transform 1 0 15088 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_162
timestamp -3600
transform 1 0 15456 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_168
timestamp -3600
transform 1 0 16008 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_176
timestamp -3600
transform 1 0 16744 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_188
timestamp -3600
transform 1 0 17848 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp -3600
transform 1 0 18676 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp -3600
transform 1 0 19044 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp -3600
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_15
timestamp -3600
transform 1 0 1932 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_19
timestamp -3600
transform 1 0 2300 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_29
timestamp -3600
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_40
timestamp -3600
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_73
timestamp -3600
transform 1 0 7268 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp -3600
transform 1 0 7636 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_129
timestamp -3600
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_159
timestamp -3600
transform 1 0 15180 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp -3600
transform 1 0 15916 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp -3600
transform 1 0 16100 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp -3600
transform 1 0 17204 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_193
timestamp -3600
transform 1 0 18308 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_201
timestamp -3600
transform 1 0 19044 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp -3600
transform 1 0 828 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp -3600
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_43
timestamp -3600
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_73
timestamp -3600
transform 1 0 7268 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_79
timestamp -3600
transform 1 0 7820 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp -3600
transform 1 0 8188 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_89
timestamp -3600
transform 1 0 8740 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_101
timestamp -3600
transform 1 0 9844 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp -3600
transform 1 0 11408 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp -3600
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_172
timestamp -3600
transform 1 0 16376 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_184
timestamp -3600
transform 1 0 17480 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp -3600
transform 1 0 18676 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp -3600
transform 1 0 19044 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp -3600
transform 1 0 828 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp -3600
transform 1 0 3036 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_39
timestamp -3600
transform 1 0 4140 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_47
timestamp -3600
transform 1 0 4876 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_52
timestamp -3600
transform 1 0 5336 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_62
timestamp -3600
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_74
timestamp -3600
transform 1 0 7360 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_90
timestamp -3600
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_94
timestamp -3600
transform 1 0 9200 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_142
timestamp -3600
transform 1 0 13616 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_191
timestamp -3600
transform 1 0 18124 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_199
timestamp -3600
transform 1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_3
timestamp -3600
transform 1 0 828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_11
timestamp -3600
transform 1 0 1564 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_18
timestamp -3600
transform 1 0 2208 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp -3600
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_29
timestamp -3600
transform 1 0 3220 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_51
timestamp -3600
transform 1 0 5244 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_55
timestamp -3600
transform 1 0 5612 0 1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp -3600
transform 1 0 6992 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp -3600
transform 1 0 8096 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp -3600
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_97
timestamp -3600
transform 1 0 9476 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_104
timestamp -3600
transform 1 0 10120 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_113
timestamp -3600
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_119
timestamp -3600
transform 1 0 11500 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_127
timestamp -3600
transform 1 0 12236 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp -3600
transform 1 0 12972 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp -3600
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp -3600
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_147
timestamp -3600
transform 1 0 14076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_155
timestamp -3600
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_179
timestamp -3600
transform 1 0 17020 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_191
timestamp -3600
transform 1 0 18124 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp -3600
transform 1 0 18492 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_197
timestamp -3600
transform 1 0 18676 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_201
timestamp -3600
transform 1 0 19044 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp -3600
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_20
timestamp -3600
transform 1 0 2392 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_32
timestamp -3600
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_36
timestamp -3600
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp -3600
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_80
timestamp -3600
transform 1 0 7912 0 -1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_92
timestamp -3600
transform 1 0 9016 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_104
timestamp -3600
transform 1 0 10120 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp -3600
transform 1 0 10948 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_119
timestamp -3600
transform 1 0 11500 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_128
timestamp -3600
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp -3600
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp -3600
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_193
timestamp -3600
transform 1 0 18308 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_201
timestamp -3600
transform 1 0 19044 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_19
timestamp -3600
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_32
timestamp -3600
transform 1 0 3496 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_43
timestamp -3600
transform 1 0 4508 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_50
timestamp -3600
transform 1 0 5152 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_78
timestamp -3600
transform 1 0 7728 0 1 14688
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_101
timestamp -3600
transform 1 0 9844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_113
timestamp -3600
transform 1 0 10948 0 1 14688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_122
timestamp -3600
transform 1 0 11776 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_134
timestamp -3600
transform 1 0 12880 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_141
timestamp -3600
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_149
timestamp -3600
transform 1 0 14260 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_163
timestamp -3600
transform 1 0 15548 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_175
timestamp -3600
transform 1 0 16652 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_187
timestamp -3600
transform 1 0 17756 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp -3600
transform 1 0 18492 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp -3600
transform 1 0 18676 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_201
timestamp -3600
transform 1 0 19044 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_36
timestamp -3600
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_48
timestamp -3600
transform 1 0 4968 0 -1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp -3600
transform 1 0 5796 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_89
timestamp -3600
transform 1 0 8740 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp -3600
transform 1 0 11684 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_132
timestamp -3600
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp -3600
transform 1 0 13156 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp -3600
transform 1 0 14260 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp -3600
transform 1 0 15364 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp -3600
transform 1 0 15916 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp -3600
transform 1 0 16100 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp -3600
transform 1 0 17204 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_193
timestamp -3600
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_201
timestamp -3600
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_3
timestamp -3600
transform 1 0 828 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_11
timestamp -3600
transform 1 0 1564 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_18
timestamp -3600
transform 1 0 2208 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp -3600
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp -3600
transform 1 0 3220 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_37
timestamp -3600
transform 1 0 3956 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp -3600
transform 1 0 4876 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_59
timestamp -3600
transform 1 0 5980 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_67
timestamp -3600
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp -3600
transform 1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_85
timestamp -3600
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_93
timestamp -3600
transform 1 0 9108 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_104
timestamp -3600
transform 1 0 10120 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_113
timestamp -3600
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_160
timestamp -3600
transform 1 0 15272 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_172
timestamp -3600
transform 1 0 16376 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_184
timestamp -3600
transform 1 0 17480 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp -3600
transform 1 0 18676 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp -3600
transform 1 0 19044 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp -3600
transform 1 0 828 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_15
timestamp -3600
transform 1 0 1932 0 -1 16864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_22
timestamp -3600
transform 1 0 2576 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_34
timestamp -3600
transform 1 0 3680 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_39
timestamp -3600
transform 1 0 4140 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_47
timestamp -3600
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_80
timestamp -3600
transform 1 0 7912 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_104
timestamp -3600
transform 1 0 10120 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp -3600
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_132
timestamp -3600
transform 1 0 12696 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_144
timestamp -3600
transform 1 0 13800 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_156
timestamp -3600
transform 1 0 14904 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp -3600
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp -3600
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_193
timestamp -3600
transform 1 0 18308 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_201
timestamp -3600
transform 1 0 19044 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp -3600
transform 1 0 828 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_11
timestamp -3600
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp -3600
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_29
timestamp -3600
transform 1 0 3220 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_37
timestamp -3600
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_46
timestamp -3600
transform 1 0 4784 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_63
timestamp -3600
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp -3600
transform 1 0 8188 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp -3600
transform 1 0 8372 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp -3600
transform 1 0 9108 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_113
timestamp -3600
transform 1 0 10948 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_125
timestamp -3600
transform 1 0 12052 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_137
timestamp -3600
transform 1 0 13156 0 1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp -3600
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp -3600
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp -3600
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp -3600
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp -3600
transform 1 0 17940 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp -3600
transform 1 0 18492 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp -3600
transform 1 0 18676 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_201
timestamp -3600
transform 1 0 19044 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_3
timestamp -3600
transform 1 0 828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_43
timestamp -3600
transform 1 0 4508 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp -3600
transform 1 0 5520 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_57
timestamp -3600
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_68
timestamp -3600
transform 1 0 6808 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_87
timestamp -3600
transform 1 0 8556 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_91
timestamp -3600
transform 1 0 8924 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_100
timestamp -3600
transform 1 0 9752 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_106
timestamp -3600
transform 1 0 10304 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp -3600
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_113
timestamp -3600
transform 1 0 10948 0 -1 17952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_121
timestamp -3600
transform 1 0 11684 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_133
timestamp -3600
transform 1 0 12788 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_145
timestamp -3600
transform 1 0 13892 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp -3600
transform 1 0 16100 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp -3600
transform 1 0 17204 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_193
timestamp -3600
transform 1 0 18308 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_201
timestamp -3600
transform 1 0 19044 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp -3600
transform 1 0 828 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp -3600
transform 1 0 1932 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp -3600
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp -3600
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_34
timestamp -3600
transform 1 0 3680 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_58
timestamp -3600
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_120
timestamp -3600
transform 1 0 11592 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_132
timestamp -3600
transform 1 0 12696 0 1 17952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp -3600
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_153
timestamp -3600
transform 1 0 14628 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_159
timestamp -3600
transform 1 0 15180 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_171
timestamp -3600
transform 1 0 16284 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp -3600
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp -3600
transform 1 0 17940 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp -3600
transform 1 0 18492 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp -3600
transform 1 0 18676 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_201
timestamp -3600
transform 1 0 19044 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp -3600
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_14
timestamp -3600
transform 1 0 1840 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_26
timestamp -3600
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_29
timestamp -3600
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_37
timestamp -3600
transform 1 0 3956 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_43
timestamp -3600
transform 1 0 4508 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp -3600
transform 1 0 5612 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_57
timestamp -3600
transform 1 0 5796 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_61
timestamp -3600
transform 1 0 6164 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_73
timestamp -3600
transform 1 0 7268 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_79
timestamp -3600
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp -3600
transform 1 0 8188 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_85
timestamp -3600
transform 1 0 8372 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_93
timestamp -3600
transform 1 0 9108 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_100
timestamp -3600
transform 1 0 9752 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_116
timestamp -3600
transform 1 0 11224 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_128
timestamp -3600
transform 1 0 12328 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_133
timestamp -3600
transform 1 0 12788 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_139
timestamp -3600
transform 1 0 13340 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_141
timestamp -3600
transform 1 0 13524 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_147
timestamp -3600
transform 1 0 14076 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_151
timestamp -3600
transform 1 0 14444 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp -3600
transform 1 0 15548 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp -3600
transform 1 0 15916 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_172
timestamp -3600
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_187
timestamp -3600
transform 1 0 17756 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_195
timestamp -3600
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_197
timestamp -3600
transform 1 0 18676 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp -3600
transform 1 0 19044 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -3600
transform -1 0 3036 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -3600
transform -1 0 3956 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -3600
transform -1 0 10948 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp -3600
transform -1 0 10212 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp -3600
transform -1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -3600
transform -1 0 16376 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -3600
transform -1 0 14444 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -3600
transform -1 0 12788 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -3600
transform 1 0 10948 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -3600
transform 1 0 9476 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -3600
transform -1 0 7820 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -3600
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp -3600
transform 1 0 4232 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input9
timestamp -3600
transform 1 0 2576 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp -3600
transform 1 0 920 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -3600
transform 1 0 17480 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap12
timestamp -3600
transform -1 0 11132 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap13
timestamp -3600
transform -1 0 10948 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap14
timestamp -3600
transform 1 0 11132 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_34
timestamp -3600
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -3600
transform -1 0 19412 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_35
timestamp -3600
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -3600
transform -1 0 19412 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_36
timestamp -3600
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -3600
transform -1 0 19412 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_37
timestamp -3600
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -3600
transform -1 0 19412 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_38
timestamp -3600
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -3600
transform -1 0 19412 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_39
timestamp -3600
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -3600
transform -1 0 19412 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_40
timestamp -3600
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -3600
transform -1 0 19412 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_41
timestamp -3600
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -3600
transform -1 0 19412 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_42
timestamp -3600
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -3600
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_43
timestamp -3600
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -3600
transform -1 0 19412 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_44
timestamp -3600
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -3600
transform -1 0 19412 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_45
timestamp -3600
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -3600
transform -1 0 19412 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_46
timestamp -3600
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -3600
transform -1 0 19412 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_47
timestamp -3600
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -3600
transform -1 0 19412 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_48
timestamp -3600
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -3600
transform -1 0 19412 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_49
timestamp -3600
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -3600
transform -1 0 19412 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_50
timestamp -3600
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -3600
transform -1 0 19412 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_51
timestamp -3600
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -3600
transform -1 0 19412 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_52
timestamp -3600
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -3600
transform -1 0 19412 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_53
timestamp -3600
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -3600
transform -1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_54
timestamp -3600
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -3600
transform -1 0 19412 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_55
timestamp -3600
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -3600
transform -1 0 19412 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_56
timestamp -3600
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -3600
transform -1 0 19412 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_57
timestamp -3600
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -3600
transform -1 0 19412 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_58
timestamp -3600
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -3600
transform -1 0 19412 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_59
timestamp -3600
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -3600
transform -1 0 19412 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_60
timestamp -3600
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -3600
transform -1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_61
timestamp -3600
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -3600
transform -1 0 19412 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_62
timestamp -3600
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -3600
transform -1 0 19412 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_63
timestamp -3600
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -3600
transform -1 0 19412 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_64
timestamp -3600
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -3600
transform -1 0 19412 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_65
timestamp -3600
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -3600
transform -1 0 19412 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_66
timestamp -3600
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp -3600
transform -1 0 19412 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_67
timestamp -3600
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp -3600
transform -1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp -3600
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp -3600
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp -3600
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp -3600
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp -3600
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp -3600
transform 1 0 16008 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_74
timestamp -3600
transform 1 0 18584 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp -3600
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp -3600
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp -3600
transform 1 0 16008 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp -3600
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp -3600
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp -3600
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp -3600
transform 1 0 18584 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp -3600
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp -3600
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp -3600
transform 1 0 16008 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_85
timestamp -3600
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp -3600
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp -3600
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp -3600
transform 1 0 18584 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_89
timestamp -3600
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_90
timestamp -3600
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp -3600
transform 1 0 16008 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_92
timestamp -3600
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_93
timestamp -3600
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_94
timestamp -3600
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp -3600
transform 1 0 18584 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_96
timestamp -3600
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_97
timestamp -3600
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_98
timestamp -3600
transform 1 0 16008 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_99
timestamp -3600
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_100
timestamp -3600
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_101
timestamp -3600
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_102
timestamp -3600
transform 1 0 18584 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_103
timestamp -3600
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_104
timestamp -3600
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_105
timestamp -3600
transform 1 0 16008 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_106
timestamp -3600
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_107
timestamp -3600
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_108
timestamp -3600
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_109
timestamp -3600
transform 1 0 18584 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_110
timestamp -3600
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_111
timestamp -3600
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_112
timestamp -3600
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_113
timestamp -3600
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_114
timestamp -3600
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_115
timestamp -3600
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_116
timestamp -3600
transform 1 0 18584 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_117
timestamp -3600
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_118
timestamp -3600
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_119
timestamp -3600
transform 1 0 16008 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_120
timestamp -3600
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_121
timestamp -3600
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_122
timestamp -3600
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_123
timestamp -3600
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_124
timestamp -3600
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_125
timestamp -3600
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_126
timestamp -3600
transform 1 0 16008 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_127
timestamp -3600
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_128
timestamp -3600
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_129
timestamp -3600
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_130
timestamp -3600
transform 1 0 18584 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_131
timestamp -3600
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_132
timestamp -3600
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_133
timestamp -3600
transform 1 0 16008 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_134
timestamp -3600
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_135
timestamp -3600
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_136
timestamp -3600
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_137
timestamp -3600
transform 1 0 18584 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_138
timestamp -3600
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_139
timestamp -3600
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_140
timestamp -3600
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_141
timestamp -3600
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_142
timestamp -3600
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_143
timestamp -3600
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_144
timestamp -3600
transform 1 0 18584 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_145
timestamp -3600
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_146
timestamp -3600
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_147
timestamp -3600
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_148
timestamp -3600
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_149
timestamp -3600
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_150
timestamp -3600
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_151
timestamp -3600
transform 1 0 18584 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_152
timestamp -3600
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_153
timestamp -3600
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_154
timestamp -3600
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_155
timestamp -3600
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_156
timestamp -3600
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_157
timestamp -3600
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_158
timestamp -3600
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_159
timestamp -3600
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_160
timestamp -3600
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_161
timestamp -3600
transform 1 0 16008 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_162
timestamp -3600
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_163
timestamp -3600
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_164
timestamp -3600
transform 1 0 13432 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_165
timestamp -3600
transform 1 0 18584 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_166
timestamp -3600
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_167
timestamp -3600
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_168
timestamp -3600
transform 1 0 16008 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_169
timestamp -3600
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_170
timestamp -3600
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_171
timestamp -3600
transform 1 0 13432 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_172
timestamp -3600
transform 1 0 18584 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_173
timestamp -3600
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_174
timestamp -3600
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_175
timestamp -3600
transform 1 0 16008 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_176
timestamp -3600
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_177
timestamp -3600
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_178
timestamp -3600
transform 1 0 13432 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_179
timestamp -3600
transform 1 0 18584 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_180
timestamp -3600
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_181
timestamp -3600
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_182
timestamp -3600
transform 1 0 16008 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_183
timestamp -3600
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_184
timestamp -3600
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_185
timestamp -3600
transform 1 0 13432 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_186
timestamp -3600
transform 1 0 18584 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_187
timestamp -3600
transform 1 0 3128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_188
timestamp -3600
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_189
timestamp -3600
transform 1 0 8280 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_190
timestamp -3600
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_191
timestamp -3600
transform 1 0 13432 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_192
timestamp -3600
transform 1 0 16008 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_193
timestamp -3600
transform 1 0 18584 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire1
timestamp -3600
transform 1 0 6440 0 -1 16864
box -38 -48 314 592
<< labels >>
rlabel metal2 s 10061 19040 10061 19040 4 VGND
rlabel metal1 s 9982 18496 9982 18496 4 VPWR
rlabel metal2 s 16698 17918 16698 17918 4 _000_
rlabel metal2 s 3353 17714 3353 17714 4 _001_
rlabel metal2 s 2346 17238 2346 17238 4 _002_
rlabel metal1 s 1145 14926 1145 14926 4 _003_
rlabel metal1 s 3496 15130 3496 15130 4 _004_
rlabel metal1 s 4564 13838 4564 13838 4 _005_
rlabel metal2 s 5566 14246 5566 14246 4 _006_
rlabel metal1 s 7084 12614 7084 12614 4 _007_
rlabel metal2 s 6670 11458 6670 11458 4 _008_
rlabel metal1 s 3905 11594 3905 11594 4 _009_
rlabel metal1 s 1973 10574 1973 10574 4 _010_
rlabel metal1 s 2157 12682 2157 12682 4 _011_
rlabel metal2 s 1329 13430 1329 13430 4 _012_
rlabel metal1 s 8142 7310 8142 7310 4 _013_
rlabel metal2 s 9618 6154 9618 6154 4 _014_
rlabel metal2 s 7682 9146 7682 9146 4 _015_
rlabel metal1 s 9250 8330 9250 8330 4 _016_
rlabel metal1 s 9885 5746 9885 5746 4 _017_
rlabel metal1 s 11352 5134 11352 5134 4 _018_
rlabel metal1 s 11403 5746 11403 5746 4 _019_
rlabel metal1 s 13662 9418 13662 9418 4 _020_
rlabel metal1 s 11990 15946 11990 15946 4 _021_
rlabel metal1 s 13478 15674 13478 15674 4 _022_
rlabel metal1 s 12834 14042 12834 14042 4 _023_
rlabel metal1 s 12036 13430 12036 13430 4 _024_
rlabel metal2 s 9982 13158 9982 13158 4 _025_
rlabel metal2 s 8510 11764 8510 11764 4 _026_
rlabel metal1 s 10994 11866 10994 11866 4 _027_
rlabel metal1 s 8873 10574 8873 10574 4 _028_
rlabel metal2 s 7866 16898 7866 16898 4 _029_
rlabel metal1 s 9966 18122 9966 18122 4 _030_
rlabel metal1 s 6711 14926 6711 14926 4 _031_
rlabel metal2 s 9425 15606 9425 15606 4 _032_
rlabel metal1 s 8157 18122 8157 18122 4 _033_
rlabel metal1 s 9752 16762 9752 16762 4 _034_
rlabel metal1 s 5857 18122 5857 18122 4 _035_
rlabel metal2 s 8970 14722 8970 14722 4 _036_
rlabel metal1 s 2514 17034 2514 17034 4 _037_
rlabel metal2 s 2530 16796 2530 16796 4 _038_
rlabel metal1 s 2116 15470 2116 15470 4 _039_
rlabel metal2 s 1334 15606 1334 15606 4 _040_
rlabel metal1 s 1012 15538 1012 15538 4 _041_
rlabel metal1 s 2530 14892 2530 14892 4 _042_
rlabel metal1 s 3082 15130 3082 15130 4 _043_
rlabel metal1 s 3174 14926 3174 14926 4 _044_
rlabel metal1 s 4600 14858 4600 14858 4 _045_
rlabel metal2 s 4186 14518 4186 14518 4 _046_
rlabel metal1 s 4830 14518 4830 14518 4 _047_
rlabel metal1 s 4692 12682 4692 12682 4 _048_
rlabel metal1 s 5152 14246 5152 14246 4 _049_
rlabel metal2 s 5382 14042 5382 14042 4 _050_
rlabel metal1 s 6164 13158 6164 13158 4 _051_
rlabel metal1 s 5290 12614 5290 12614 4 _052_
rlabel metal1 s 5980 12138 5980 12138 4 _053_
rlabel metal1 s 5336 11866 5336 11866 4 _054_
rlabel metal1 s 5398 11594 5398 11594 4 _055_
rlabel metal1 s 5980 11186 5980 11186 4 _056_
rlabel metal1 s 2530 11628 2530 11628 4 _057_
rlabel metal2 s 4094 11696 4094 11696 4 _058_
rlabel metal2 s 4278 11798 4278 11798 4 _059_
rlabel metal2 s 3174 11968 3174 11968 4 _060_
rlabel metal1 s 2576 11254 2576 11254 4 _061_
rlabel metal1 s 2116 11186 2116 11186 4 _062_
rlabel metal1 s 2300 13362 2300 13362 4 _063_
rlabel metal2 s 2898 12580 2898 12580 4 _064_
rlabel metal1 s 1886 13872 1886 13872 4 _065_
rlabel metal1 s 8418 7174 8418 7174 4 _066_
rlabel metal2 s 9522 9452 9522 9452 4 _067_
rlabel metal2 s 9982 9792 9982 9792 4 _068_
rlabel metal1 s 9338 9486 9338 9486 4 _069_
rlabel metal1 s 16560 13362 16560 13362 4 _070_
rlabel metal1 s 11270 9554 11270 9554 4 _071_
rlabel metal1 s 15502 8398 15502 8398 4 _072_
rlabel metal1 s 14858 11152 14858 11152 4 _073_
rlabel metal1 s 17296 9146 17296 9146 4 _074_
rlabel metal1 s 17158 10438 17158 10438 4 _075_
rlabel metal1 s 15226 13192 15226 13192 4 _076_
rlabel metal2 s 18354 8806 18354 8806 4 _077_
rlabel metal1 s 15364 11662 15364 11662 4 _078_
rlabel metal1 s 17411 8398 17411 8398 4 _079_
rlabel metal1 s 16100 11866 16100 11866 4 _080_
rlabel metal2 s 14122 7786 14122 7786 4 _081_
rlabel metal1 s 16956 8398 16956 8398 4 _082_
rlabel metal2 s 13478 11254 13478 11254 4 _083_
rlabel metal1 s 16790 8432 16790 8432 4 _084_
rlabel metal1 s 15226 8500 15226 8500 4 _085_
rlabel metal1 s 13708 11186 13708 11186 4 _086_
rlabel metal1 s 15870 8364 15870 8364 4 _087_
rlabel metal1 s 15686 8058 15686 8058 4 _088_
rlabel metal2 s 16054 7582 16054 7582 4 _089_
rlabel metal1 s 12512 8398 12512 8398 4 _090_
rlabel metal1 s 15134 8364 15134 8364 4 _091_
rlabel metal2 s 17342 9010 17342 9010 4 _092_
rlabel metal1 s 16008 9146 16008 9146 4 _093_
rlabel metal1 s 16054 8058 16054 8058 4 _094_
rlabel metal2 s 15410 8636 15410 8636 4 _095_
rlabel metal2 s 14950 8024 14950 8024 4 _096_
rlabel metal1 s 8464 7310 8464 7310 4 _097_
rlabel metal1 s 11914 16628 11914 16628 4 _098_
rlabel metal2 s 12006 13906 12006 13906 4 _099_
rlabel metal1 s 8970 18598 8970 18598 4 _100_
rlabel metal2 s 13754 9248 13754 9248 4 _101_
rlabel metal2 s 15502 12988 15502 12988 4 _102_
rlabel metal1 s 16100 10166 16100 10166 4 _103_
rlabel metal2 s 16330 9690 16330 9690 4 _104_
rlabel metal2 s 15318 8092 15318 8092 4 _105_
rlabel metal2 s 16422 6970 16422 6970 4 _106_
rlabel metal2 s 15226 6766 15226 6766 4 _107_
rlabel metal1 s 16606 11152 16606 11152 4 _108_
rlabel metal2 s 16882 11356 16882 11356 4 _109_
rlabel metal1 s 14674 10574 14674 10574 4 _110_
rlabel metal2 s 15571 6902 15571 6902 4 _111_
rlabel metal1 s 14398 6800 14398 6800 4 _112_
rlabel metal2 s 14306 7140 14306 7140 4 _113_
rlabel metal1 s 15134 6766 15134 6766 4 _114_
rlabel metal1 s 14122 6664 14122 6664 4 _115_
rlabel metal1 s 8832 6834 8832 6834 4 _116_
rlabel metal1 s 7452 9146 7452 9146 4 _117_
rlabel metal2 s 13202 9826 13202 9826 4 _118_
rlabel metal1 s 14674 11220 14674 11220 4 _119_
rlabel metal1 s 13938 11050 13938 11050 4 _120_
rlabel metal2 s 14490 10880 14490 10880 4 _121_
rlabel metal2 s 13294 10438 13294 10438 4 _122_
rlabel metal2 s 15134 10778 15134 10778 4 _123_
rlabel metal1 s 13386 10132 13386 10132 4 _124_
rlabel metal1 s 14260 10166 14260 10166 4 _125_
rlabel metal1 s 14214 8364 14214 8364 4 _126_
rlabel metal1 s 13524 8466 13524 8466 4 _127_
rlabel metal2 s 13662 10047 13662 10047 4 _128_
rlabel metal1 s 14260 9690 14260 9690 4 _129_
rlabel metal1 s 13616 10030 13616 10030 4 _130_
rlabel metal2 s 13018 9758 13018 9758 4 _131_
rlabel metal1 s 7452 9010 7452 9010 4 _132_
rlabel metal1 s 13478 8058 13478 8058 4 _133_
rlabel metal2 s 13570 7378 13570 7378 4 _134_
rlabel metal1 s 13202 7888 13202 7888 4 _135_
rlabel metal1 s 12880 8058 12880 8058 4 _136_
rlabel metal1 s 12052 8602 12052 8602 4 _137_
rlabel metal2 s 11914 9180 11914 9180 4 _138_
rlabel metal1 s 10534 8976 10534 8976 4 _139_
rlabel metal1 s 17710 8942 17710 8942 4 _140_
rlabel metal1 s 14720 9078 14720 9078 4 _141_
rlabel metal1 s 13248 8602 13248 8602 4 _142_
rlabel metal1 s 12512 8806 12512 8806 4 _143_
rlabel metal1 s 10350 9044 10350 9044 4 _144_
rlabel metal1 s 9660 9146 9660 9146 4 _145_
rlabel metal1 s 9844 16014 9844 16014 4 _146_
rlabel metal1 s 9246 9010 9246 9010 4 _147_
rlabel metal1 s 9568 17510 9568 17510 4 _148_
rlabel metal1 s 12190 6970 12190 6970 4 _149_
rlabel metal1 s 13202 7242 13202 7242 4 _150_
rlabel metal1 s 10672 7446 10672 7446 4 _151_
rlabel metal1 s 13570 7310 13570 7310 4 _152_
rlabel metal1 s 12742 7208 12742 7208 4 _153_
rlabel metal1 s 11178 6766 11178 6766 4 _154_
rlabel metal2 s 9982 6426 9982 6426 4 _155_
rlabel metal3 s 10189 16660 10189 16660 4 _156_
rlabel metal1 s 13018 6970 13018 6970 4 _157_
rlabel metal1 s 10994 7378 10994 7378 4 _158_
rlabel metal2 s 11040 6834 11040 6834 4 _159_
rlabel metal1 s 10580 6222 10580 6222 4 _160_
rlabel metal2 s 10350 6698 10350 6698 4 _161_
rlabel metal1 s 10672 15334 10672 15334 4 _162_
rlabel metal2 s 11638 16218 11638 16218 4 _163_
rlabel metal2 s 11546 15946 11546 15946 4 _164_
rlabel metal1 s 11746 14858 11746 14858 4 _165_
rlabel metal2 s 12926 15334 12926 15334 4 _166_
rlabel metal1 s 12466 13940 12466 13940 4 _167_
rlabel metal1 s 12788 13838 12788 13838 4 _168_
rlabel metal1 s 12696 12410 12696 12410 4 _169_
rlabel metal2 s 11822 13532 11822 13532 4 _170_
rlabel metal2 s 11730 13124 11730 13124 4 _171_
rlabel metal1 s 11178 12954 11178 12954 4 _172_
rlabel metal1 s 10948 13838 10948 13838 4 _173_
rlabel metal1 s 10212 12750 10212 12750 4 _174_
rlabel metal1 s 9108 12886 9108 12886 4 _175_
rlabel metal1 s 10764 12886 10764 12886 4 _176_
rlabel metal2 s 10902 11866 10902 11866 4 _177_
rlabel metal1 s 9752 10982 9752 10982 4 _178_
rlabel metal1 s 10074 11050 10074 11050 4 _179_
rlabel metal1 s 9430 11186 9430 11186 4 _180_
rlabel metal1 s 7590 18190 7590 18190 4 _181_
rlabel metal1 s 7176 16762 7176 16762 4 _182_
rlabel metal2 s 9062 18088 9062 18088 4 _183_
rlabel metal2 s 7866 15232 7866 15232 4 _184_
rlabel metal1 s 9430 16048 9430 16048 4 _185_
rlabel metal1 s 8464 17850 8464 17850 4 _186_
rlabel metal1 s 9108 16762 9108 16762 4 _187_
rlabel metal1 s 6486 17850 6486 17850 4 _188_
rlabel metal1 s 8418 14586 8418 14586 4 _189_
rlabel metal1 s 3910 17238 3910 17238 4 _190_
rlabel metal1 s 8234 13362 8234 13362 4 _191_
rlabel metal2 s 8326 13124 8326 13124 4 _192_
rlabel metal2 s 4462 13090 4462 13090 4 _193_
rlabel metal1 s 7222 13362 7222 13362 4 _194_
rlabel metal1 s 10994 15436 10994 15436 4 _195_
rlabel metal1 s 5060 16218 5060 16218 4 _196_
rlabel metal1 s 6072 17306 6072 17306 4 _197_
rlabel metal2 s 9338 17952 9338 17952 4 _198_
rlabel metal1 s 4922 17136 4922 17136 4 _199_
rlabel metal1 s 5474 16626 5474 16626 4 _200_
rlabel metal2 s 8878 16864 8878 16864 4 _201_
rlabel metal2 s 5658 17306 5658 17306 4 _202_
rlabel metal1 s 5566 16558 5566 16558 4 _203_
rlabel metal1 s 5198 16660 5198 16660 4 _204_
rlabel metal1 s 6486 16558 6486 16558 4 _205_
rlabel metal2 s 11362 15844 11362 15844 4 _206_
rlabel metal1 s 8372 14518 8372 14518 4 _207_
rlabel metal2 s 2622 15215 2622 15215 4 _208_
rlabel metal1 s 3588 17306 3588 17306 4 _209_
rlabel metal1 s 2576 17306 2576 17306 4 _210_
rlabel metal3 s 18515 15980 18515 15980 4 clk
rlabel metal3 s 10580 12716 10580 12716 4 clknet_0_clk
rlabel metal1 s 1932 12750 1932 12750 4 clknet_2_0__leaf_clk
rlabel metal1 s 1242 17646 1242 17646 4 clknet_2_1__leaf_clk
rlabel metal1 s 14605 5746 14605 5746 4 clknet_2_2__leaf_clk
rlabel metal2 s 13570 16864 13570 16864 4 clknet_2_3__leaf_clk
rlabel metal1 s 16054 18802 16054 18802 4 data[0]
rlabel metal1 s 14260 18802 14260 18802 4 data[1]
rlabel metal1 s 12604 18802 12604 18802 4 data[2]
rlabel metal1 s 10994 18802 10994 18802 4 data[3]
rlabel metal1 s 9706 18836 9706 18836 4 data[4]
rlabel metal1 s 7544 18802 7544 18802 4 data[5]
rlabel metal1 s 5888 18802 5888 18802 4 data[6]
rlabel metal1 s 4232 18802 4232 18802 4 data[7]
rlabel metal1 s 2576 18802 2576 18802 4 ext_data
rlabel metal1 s 920 18802 920 18802 4 load_divider
rlabel metal1 s 17572 18802 17572 18802 4 n_rst
rlabel metal1 s 14306 17612 14306 17612 4 net1
rlabel metal2 s 6486 18190 6486 18190 4 net10
rlabel metal2 s 16790 18394 16790 18394 4 net11
rlabel metal1 s 10626 12750 10626 12750 4 net12
rlabel metal2 s 8878 11390 8878 11390 4 net13
rlabel metal1 s 11638 16524 11638 16524 4 net14
rlabel metal2 s 14490 17918 14490 17918 4 net15
rlabel metal2 s 2346 13600 2346 13600 4 net16
rlabel metal1 s 3220 12614 3220 12614 4 net17
rlabel metal1 s 10120 15878 10120 15878 4 net18
rlabel metal1 s 8970 11220 8970 11220 4 net19
rlabel metal1 s 13317 18666 13317 18666 4 net2
rlabel metal1 s 10718 12818 10718 12818 4 net20
rlabel metal1 s 11178 16694 11178 16694 4 net21
rlabel metal2 s 12558 17408 12558 17408 4 net3
rlabel metal2 s 10626 18156 10626 18156 4 net4
rlabel metal2 s 9522 18156 9522 18156 4 net5
rlabel metal1 s 9430 16626 9430 16626 4 net6
rlabel metal1 s 6670 18258 6670 18258 4 net7
rlabel metal1 s 8694 14348 8694 14348 4 net8
rlabel metal1 s 8464 18802 8464 18802 4 net9
rlabel metal2 s 1242 1928 1242 1928 4 r2r_out[0]
rlabel metal1 s 6118 4114 6118 4114 4 r2r_out[1]
rlabel metal1 s 6394 9350 6394 9350 4 r2r_out[2]
rlabel metal1 s 8602 8534 8602 8534 4 r2r_out[3]
rlabel metal1 s 10948 5542 10948 5542 4 r2r_out[4]
rlabel metal1 s 13110 4998 13110 4998 4 r2r_out[5]
rlabel metal2 s 16146 2948 16146 2948 4 r2r_out[6]
rlabel metal1 s 18400 5542 18400 5542 4 r2r_out[7]
rlabel metal1 s 2208 17102 2208 17102 4 sine_lookup.count\[0\]
rlabel metal1 s 2668 12614 2668 12614 4 sine_lookup.count\[10\]
rlabel metal2 s 4002 12920 4002 12920 4 sine_lookup.count\[11\]
rlabel metal2 s 5014 17102 5014 17102 4 sine_lookup.count\[1\]
rlabel metal1 s 2200 14518 2200 14518 4 sine_lookup.count\[2\]
rlabel metal2 s 2438 15844 2438 15844 4 sine_lookup.count\[3\]
rlabel metal1 s 4140 14926 4140 14926 4 sine_lookup.count\[4\]
rlabel metal2 s 6118 16643 6118 16643 4 sine_lookup.count\[5\]
rlabel metal1 s 5290 13294 5290 13294 4 sine_lookup.count\[6\]
rlabel metal1 s 8234 13430 8234 13430 4 sine_lookup.count\[7\]
rlabel metal2 s 4922 12410 4922 12410 4 sine_lookup.count\[8\]
rlabel metal1 s 3404 12954 3404 12954 4 sine_lookup.count\[9\]
rlabel metal1 s 6716 17102 6716 17102 4 sine_lookup.divider\[0\]
rlabel metal1 s 11316 18190 11316 18190 4 sine_lookup.divider\[1\]
rlabel metal2 s 7314 14212 7314 14212 4 sine_lookup.divider\[2\]
rlabel metal1 s 10810 16150 10810 16150 4 sine_lookup.divider\[3\]
rlabel metal2 s 6854 17646 6854 17646 4 sine_lookup.divider\[4\]
rlabel metal1 s 10672 17102 10672 17102 4 sine_lookup.divider\[5\]
rlabel metal2 s 5014 17850 5014 17850 4 sine_lookup.divider\[6\]
rlabel metal1 s 8740 15130 8740 15130 4 sine_lookup.divider\[7\]
rlabel metal1 s 14191 17850 14191 17850 4 sine_lookup.rst
rlabel metal2 s 14950 14688 14950 14688 4 sine_lookup.sine_input\[0\]
rlabel metal2 s 16238 13600 16238 13600 4 sine_lookup.sine_input\[1\]
rlabel metal2 s 15134 13056 15134 13056 4 sine_lookup.sine_input\[2\]
rlabel metal1 s 13616 13158 13616 13158 4 sine_lookup.sine_input\[3\]
rlabel metal1 s 11546 13260 11546 13260 4 sine_lookup.sine_input\[4\]
rlabel metal2 s 8326 11458 8326 11458 4 sine_lookup.sine_input\[5\]
rlabel metal1 s 14122 12206 14122 12206 4 sine_lookup.sine_input\[6\]
rlabel metal1 s 10166 10166 10166 10166 4 sine_lookup.sine_input\[7\]
flabel metal4 s 19251 496 19571 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 14536 496 14856 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 9821 496 10141 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5106 496 5426 19088 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 16894 496 17214 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 12179 496 12499 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7464 496 7784 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2749 496 3069 19088 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 19062 19600 19118 20000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 15750 19600 15806 20000 0 FreeSans 280 90 0 0 data[0]
port 4 nsew
flabel metal2 s 14094 19600 14150 20000 0 FreeSans 280 90 0 0 data[1]
port 5 nsew
flabel metal2 s 12438 19600 12494 20000 0 FreeSans 280 90 0 0 data[2]
port 6 nsew
flabel metal2 s 10782 19600 10838 20000 0 FreeSans 280 90 0 0 data[3]
port 7 nsew
flabel metal2 s 9126 19600 9182 20000 0 FreeSans 280 90 0 0 data[4]
port 8 nsew
flabel metal2 s 7470 19600 7526 20000 0 FreeSans 280 90 0 0 data[5]
port 9 nsew
flabel metal2 s 5814 19600 5870 20000 0 FreeSans 280 90 0 0 data[6]
port 10 nsew
flabel metal2 s 4158 19600 4214 20000 0 FreeSans 280 90 0 0 data[7]
port 11 nsew
flabel metal2 s 2502 19600 2558 20000 0 FreeSans 280 90 0 0 ext_data
port 12 nsew
flabel metal2 s 846 19600 902 20000 0 FreeSans 280 90 0 0 load_divider
port 13 nsew
flabel metal2 s 17406 19600 17462 20000 0 FreeSans 280 90 0 0 n_rst
port 14 nsew
flabel metal2 s 1214 0 1270 400 0 FreeSans 280 90 0 0 r2r_out[0]
port 15 nsew
flabel metal2 s 3698 0 3754 400 0 FreeSans 280 90 0 0 r2r_out[1]
port 16 nsew
flabel metal2 s 6182 0 6238 400 0 FreeSans 280 90 0 0 r2r_out[2]
port 17 nsew
flabel metal2 s 8666 0 8722 400 0 FreeSans 280 90 0 0 r2r_out[3]
port 18 nsew
flabel metal2 s 11150 0 11206 400 0 FreeSans 280 90 0 0 r2r_out[4]
port 19 nsew
flabel metal2 s 13634 0 13690 400 0 FreeSans 280 90 0 0 r2r_out[5]
port 20 nsew
flabel metal2 s 16118 0 16174 400 0 FreeSans 280 90 0 0 r2r_out[6]
port 21 nsew
flabel metal2 s 18602 0 18658 400 0 FreeSans 280 90 0 0 r2r_out[7]
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string GDS_END 1210514
string GDS_FILE ../gds/r2r_dac_control.gds
string GDS_START 451048
<< end >>
