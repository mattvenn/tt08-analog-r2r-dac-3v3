magic
tech sky130A
magscale 1 2
timestamp 1720524744
<< metal1 >>
rect 5624 20526 5630 20738
rect 5842 20526 5848 20738
rect 8424 20526 8430 20738
rect 8642 20526 8648 20738
rect 11224 20526 11230 20738
rect 11442 20526 11448 20738
rect 14024 20526 14030 20738
rect 14242 20526 14248 20738
rect 16824 20526 16830 20738
rect 17042 20526 17048 20738
rect 19624 20526 19630 20738
rect 19842 20526 19848 20738
rect 22424 20526 22430 20738
rect 22642 20526 22648 20738
rect 25224 20526 25230 20738
rect 25442 20526 25448 20738
rect 5066 20372 5072 20428
rect 5128 20372 5134 20428
rect 4314 19946 4320 20158
rect 4532 19946 4538 20158
rect 4320 19058 4532 19946
rect 5072 19272 5128 20372
rect 5630 19158 5842 20526
rect 7866 20372 7872 20428
rect 7928 20372 7934 20428
rect 7114 19946 7120 20158
rect 7332 19946 7338 20158
rect 6227 19019 6233 19210
rect 6424 19019 6430 19210
rect 7120 19058 7332 19946
rect 7872 19172 7928 20372
rect 8430 19158 8642 20526
rect 10691 20353 10697 20409
rect 10753 20353 10759 20409
rect 9914 19946 9920 20158
rect 10132 19946 10138 20158
rect 9027 19019 9033 19210
rect 9224 19019 9230 19210
rect 9920 19058 10132 19946
rect 10697 19217 10753 20353
rect 11230 19158 11442 20526
rect 13469 20342 13475 20398
rect 13531 20342 13537 20398
rect 12714 19946 12720 20158
rect 12932 19946 12938 20158
rect 11827 19019 11833 19210
rect 12024 19019 12030 19210
rect 12720 19058 12932 19946
rect 13475 19286 13531 20342
rect 14030 19158 14242 20526
rect 16258 20365 16264 20421
rect 16320 20365 16326 20421
rect 15514 19946 15520 20158
rect 15732 19946 15738 20158
rect 14627 19019 14633 19210
rect 14824 19019 14830 19210
rect 15520 19058 15732 19946
rect 16264 19263 16320 20365
rect 16830 19158 17042 20526
rect 19082 20376 19088 20432
rect 19144 20376 19150 20432
rect 18314 19946 18320 20158
rect 18532 19946 18538 20158
rect 17427 19019 17433 19210
rect 17624 19019 17630 19210
rect 18320 19058 18532 19946
rect 19088 19217 19144 20376
rect 19630 19158 19842 20526
rect 21912 20432 21968 20438
rect 21114 19946 21120 20158
rect 21332 19946 21338 20158
rect 20227 19019 20233 19210
rect 20424 19019 20430 19210
rect 21120 19058 21332 19946
rect 21912 19251 21968 20376
rect 22430 19158 22642 20526
rect 24720 20356 24726 20412
rect 24782 20356 24788 20412
rect 23914 19946 23920 20158
rect 24132 19946 24138 20158
rect 23027 19019 23033 19210
rect 23224 19019 23230 19210
rect 23920 19058 24132 19946
rect 24726 19232 24782 20356
rect 25230 19158 25442 20526
rect 25827 19019 25833 19210
rect 26024 19019 26030 19210
rect 6233 18787 6424 19019
rect 9033 18787 9224 19019
rect 11833 18787 12024 19019
rect 14633 18787 14824 19019
rect 17433 18787 17624 19019
rect 20233 18787 20424 19019
rect 23033 18787 23224 19019
rect 25833 18787 26024 19019
rect 5158 13066 5458 15202
rect 7978 13562 8278 15096
rect 10776 14092 11076 15202
rect 10776 13792 13464 14092
rect 7978 13262 11964 13562
rect 5158 12766 8964 13066
rect 8664 12168 8964 12766
rect 11664 12168 11964 13262
rect 13164 12168 13464 13792
rect 13928 13526 14228 15272
rect 13928 13226 14964 13526
rect 14664 12168 14964 13226
rect 16164 12164 16464 15190
rect 19098 14446 19398 15142
rect 17664 14146 19398 14446
rect 17664 12168 17964 14146
rect 21942 13750 22242 15108
rect 19164 13450 22242 13750
rect 19164 12168 19464 13450
rect 19964 13042 20264 13048
rect 24822 12970 25122 15202
rect 19964 12168 20264 12742
rect 20664 12670 25122 12970
rect 20664 12168 20964 12670
rect 5462 2520 5862 2526
rect 5862 2120 7872 2520
rect 5462 2114 5862 2120
<< via1 >>
rect 5630 20526 5842 20738
rect 8430 20526 8642 20738
rect 11230 20526 11442 20738
rect 14030 20526 14242 20738
rect 16830 20526 17042 20738
rect 19630 20526 19842 20738
rect 22430 20526 22642 20738
rect 25230 20526 25442 20738
rect 5072 20372 5128 20428
rect 4320 19946 4532 20158
rect 7872 20372 7928 20428
rect 7120 19946 7332 20158
rect 6233 19019 6424 19210
rect 10697 20353 10753 20409
rect 9920 19946 10132 20158
rect 9033 19019 9224 19210
rect 13475 20342 13531 20398
rect 12720 19946 12932 20158
rect 11833 19019 12024 19210
rect 16264 20365 16320 20421
rect 15520 19946 15732 20158
rect 14633 19019 14824 19210
rect 19088 20376 19144 20432
rect 18320 19946 18532 20158
rect 17433 19019 17624 19210
rect 21912 20376 21968 20432
rect 21120 19946 21332 20158
rect 20233 19019 20424 19210
rect 24726 20356 24782 20412
rect 23920 19946 24132 20158
rect 23033 19019 23224 19210
rect 25833 19019 26024 19210
rect 19964 12742 20264 13042
rect 5462 2120 5862 2520
<< metal2 >>
rect 14263 44154 14319 44161
rect 9796 44152 14321 44154
rect 9796 44096 14263 44152
rect 14319 44096 14321 44152
rect 9796 44094 14321 44096
rect 8470 43669 8526 43676
rect 4287 43667 8528 43669
rect 4287 43611 8470 43667
rect 8526 43611 8528 43667
rect 4287 43609 8528 43611
rect 4287 42633 4347 43609
rect 8470 43602 8526 43609
rect 8901 43459 8957 43466
rect 5934 43457 8959 43459
rect 5934 43401 8901 43457
rect 8957 43401 8959 43457
rect 5934 43399 8959 43401
rect 5934 42704 5994 43399
rect 8901 43392 8957 43399
rect 9200 43273 9256 43280
rect 7589 43271 9258 43273
rect 7589 43215 9200 43271
rect 9256 43215 9258 43271
rect 7589 43213 9258 43215
rect 7589 42595 7649 43213
rect 9200 43206 9256 43213
rect 9796 42850 9856 44094
rect 14263 44087 14319 44094
rect 14893 43978 14949 43985
rect 9211 42790 9856 42850
rect 10901 43976 14951 43978
rect 10901 43920 14893 43976
rect 14949 43920 14951 43976
rect 10901 43918 14951 43920
rect 10901 42623 10961 43918
rect 14893 43911 14949 43918
rect 16594 43821 16650 43828
rect 12560 43819 16652 43821
rect 12560 43763 16594 43819
rect 16650 43763 16652 43819
rect 12560 43761 16652 43763
rect 12560 42652 12620 43761
rect 16594 43754 16650 43761
rect 17223 43669 17279 43676
rect 14204 43667 17281 43669
rect 14204 43611 17223 43667
rect 17279 43611 17281 43667
rect 14204 43609 17281 43611
rect 14204 42671 14264 43609
rect 17223 43602 17279 43609
rect 18461 43526 18517 43533
rect 15870 43524 18519 43526
rect 15870 43468 18461 43524
rect 18517 43468 18519 43524
rect 15870 43466 18519 43468
rect 15870 42685 15930 43466
rect 18461 43459 18517 43466
rect 18171 43340 18227 43347
rect 17526 43338 18229 43340
rect 17526 43282 18171 43338
rect 18227 43282 18229 43338
rect 17526 43280 18229 43282
rect 17526 42652 17586 43280
rect 18171 43273 18227 43280
rect 21653 43162 21713 43164
rect 20208 43150 20264 43157
rect 19173 43148 20266 43150
rect 19173 43092 20208 43148
rect 20264 43092 20266 43148
rect 21646 43106 21655 43162
rect 21711 43106 21720 43162
rect 19173 43090 20266 43092
rect 19173 42752 19233 43090
rect 20208 43083 20264 43090
rect 21653 42750 21713 43106
rect 23558 42812 23614 42819
rect 22486 42810 23616 42812
rect 22486 42754 23558 42810
rect 23614 42754 23616 42810
rect 22486 42752 23616 42754
rect 20796 42690 21713 42750
rect 23558 42745 23614 42752
rect 4633 22928 5128 22984
rect 7136 22933 7928 22989
rect 4320 20527 4532 20532
rect 4316 20325 4325 20527
rect 4527 20325 4536 20527
rect 5072 20428 5128 22928
rect 5630 21469 5842 21474
rect 5626 21267 5635 21469
rect 5837 21267 5846 21469
rect 5630 20738 5842 21267
rect 7120 20527 7332 20532
rect 5630 20520 5842 20526
rect 5072 20366 5128 20372
rect 7116 20325 7125 20527
rect 7327 20325 7336 20527
rect 7872 20428 7928 22933
rect 9550 22914 10753 22970
rect 8430 21469 8642 21474
rect 8426 21267 8435 21469
rect 8637 21267 8646 21469
rect 8430 20738 8642 21267
rect 9920 20527 10132 20532
rect 8430 20520 8642 20526
rect 7872 20366 7928 20372
rect 9916 20325 9925 20527
rect 10127 20325 10136 20527
rect 10697 20409 10753 22914
rect 12087 22909 13531 22965
rect 14558 22909 16320 22965
rect 17033 22918 19144 22974
rect 11230 21469 11442 21474
rect 11226 21267 11235 21469
rect 11437 21267 11446 21469
rect 11230 20738 11442 21267
rect 12720 20527 12932 20532
rect 11230 20520 11442 20526
rect 10697 20347 10753 20353
rect 12716 20325 12725 20527
rect 12927 20325 12936 20527
rect 13475 20398 13531 22909
rect 14030 21469 14242 21474
rect 14026 21267 14035 21469
rect 14237 21267 14246 21469
rect 14030 20738 14242 21267
rect 15520 20527 15732 20532
rect 14030 20520 14242 20526
rect 13475 20336 13531 20342
rect 15516 20325 15525 20527
rect 15727 20325 15736 20527
rect 16264 20421 16320 22909
rect 16830 21469 17042 21474
rect 16826 21267 16835 21469
rect 17037 21267 17046 21469
rect 16830 20738 17042 21267
rect 18320 20527 18532 20532
rect 16830 20520 17042 20526
rect 16264 20359 16320 20365
rect 18316 20325 18325 20527
rect 18527 20325 18536 20527
rect 19088 20432 19144 22918
rect 19561 22360 19617 23079
rect 21973 22952 24782 23008
rect 21912 22360 21968 22373
rect 19561 22304 21968 22360
rect 19630 21469 19842 21474
rect 19626 21267 19635 21469
rect 19837 21267 19846 21469
rect 19630 20738 19842 21267
rect 21120 20527 21332 20532
rect 19630 20520 19842 20526
rect 19088 20370 19144 20376
rect 21116 20325 21125 20527
rect 21327 20325 21336 20527
rect 21912 20432 21968 22304
rect 22430 21469 22642 21474
rect 22426 21267 22435 21469
rect 22637 21267 22646 21469
rect 22430 20738 22642 21267
rect 23920 20527 24132 20532
rect 22430 20520 22642 20526
rect 21906 20376 21912 20432
rect 21968 20376 21974 20432
rect 23916 20325 23925 20527
rect 24127 20325 24136 20527
rect 24726 20412 24782 22952
rect 25230 21469 25442 21474
rect 25226 21267 25235 21469
rect 25437 21267 25446 21469
rect 25230 20738 25442 21267
rect 25230 20520 25442 20526
rect 24726 20350 24782 20356
rect 4320 20158 4532 20325
rect 4320 19940 4532 19946
rect 7120 20158 7332 20325
rect 7120 19940 7332 19946
rect 9920 20158 10132 20325
rect 9920 19940 10132 19946
rect 12720 20158 12932 20325
rect 12720 19940 12932 19946
rect 15520 20158 15732 20325
rect 15520 19940 15732 19946
rect 18320 20158 18532 20325
rect 18320 19940 18532 19946
rect 21120 20158 21332 20325
rect 21120 19940 21332 19946
rect 23920 20158 24132 20325
rect 23920 19940 24132 19946
rect 6233 19521 6424 19526
rect 9033 19521 9224 19526
rect 11833 19521 12024 19526
rect 14633 19521 14824 19526
rect 17433 19521 17624 19526
rect 20233 19521 20424 19526
rect 23033 19521 23224 19526
rect 25833 19521 26024 19526
rect 6229 19340 6238 19521
rect 6419 19340 6428 19521
rect 9029 19340 9038 19521
rect 9219 19340 9228 19521
rect 11829 19340 11838 19521
rect 12019 19340 12028 19521
rect 14629 19340 14638 19521
rect 14819 19340 14828 19521
rect 17429 19340 17438 19521
rect 17619 19340 17628 19521
rect 20229 19340 20238 19521
rect 20419 19340 20428 19521
rect 23029 19340 23038 19521
rect 23219 19340 23228 19521
rect 25829 19340 25838 19521
rect 26019 19340 26028 19521
rect 6233 19210 6424 19340
rect 6233 19013 6424 19019
rect 9033 19210 9224 19340
rect 9033 19013 9224 19019
rect 11833 19210 12024 19340
rect 11833 19013 12024 19019
rect 14633 19210 14824 19340
rect 14633 19013 14824 19019
rect 17433 19210 17624 19340
rect 17433 19013 17624 19019
rect 20233 19210 20424 19340
rect 20233 19013 20424 19019
rect 23033 19210 23224 19340
rect 23033 19013 23224 19019
rect 25833 19210 26024 19340
rect 25833 19013 26024 19019
rect 19958 12742 19964 13042
rect 20264 12742 23222 13042
rect 4966 10936 8488 11336
rect 4966 2524 5366 10936
rect 4569 2520 5366 2524
rect 4564 2515 5462 2520
rect 4564 2125 4569 2515
rect 4959 2125 5462 2515
rect 4564 2120 5462 2125
rect 5862 2120 5868 2520
rect 22925 2240 23220 12742
rect 4569 2116 4959 2120
rect 22925 1945 27174 2240
rect 27469 1945 27478 2240
<< via2 >>
rect 14263 44096 14319 44152
rect 8470 43611 8526 43667
rect 8901 43401 8957 43457
rect 9200 43215 9256 43271
rect 14893 43920 14949 43976
rect 16594 43763 16650 43819
rect 17223 43611 17279 43667
rect 18461 43468 18517 43524
rect 18171 43282 18227 43338
rect 20208 43092 20264 43148
rect 21655 43106 21711 43162
rect 23558 42754 23614 42810
rect 4325 20325 4527 20527
rect 5635 21267 5837 21469
rect 7125 20325 7327 20527
rect 8435 21267 8637 21469
rect 9925 20325 10127 20527
rect 11235 21267 11437 21469
rect 12725 20325 12927 20527
rect 14035 21267 14237 21469
rect 15525 20325 15727 20527
rect 16835 21267 17037 21469
rect 18325 20325 18527 20527
rect 19635 21267 19837 21469
rect 21125 20325 21327 20527
rect 22435 21267 22637 21469
rect 23925 20325 24127 20527
rect 25235 21267 25437 21469
rect 6238 19340 6419 19521
rect 9038 19340 9219 19521
rect 11838 19340 12019 19521
rect 14638 19340 14819 19521
rect 17438 19340 17619 19521
rect 20238 19340 20419 19521
rect 23038 19340 23219 19521
rect 25838 19340 26019 19521
rect 4569 2125 4959 2515
rect 27174 1945 27469 2240
<< metal3 >>
rect 16654 44794 16718 44800
rect 16718 44732 26008 44792
rect 16654 44724 16718 44730
rect 8466 44632 8530 44638
rect 8466 44562 8530 44568
rect 8468 43672 8528 44562
rect 14189 44494 14253 44500
rect 8899 44432 14189 44492
rect 8465 43667 8531 43672
rect 8465 43611 8470 43667
rect 8526 43611 8531 43667
rect 8465 43606 8531 43611
rect 8899 43462 8959 44432
rect 14189 44424 14253 44430
rect 14236 44346 14300 44352
rect 9198 44284 14236 44344
rect 8896 43457 8962 43462
rect 8896 43401 8901 43457
rect 8957 43401 8962 43457
rect 8896 43396 8962 43401
rect 9198 43276 9258 44284
rect 14236 44276 14300 44282
rect 14258 44154 14324 44157
rect 19514 44156 19578 44162
rect 14258 44152 19514 44154
rect 14258 44096 14263 44152
rect 14319 44096 19514 44152
rect 14258 44094 19514 44096
rect 14258 44091 14324 44094
rect 19514 44086 19578 44092
rect 14888 43978 14954 43981
rect 19706 43980 19770 43986
rect 14888 43976 19706 43978
rect 14888 43920 14893 43976
rect 14949 43920 19706 43976
rect 14888 43918 19706 43920
rect 14888 43915 14954 43918
rect 19706 43910 19770 43916
rect 16589 43821 16655 43824
rect 19903 43823 19967 43829
rect 16589 43819 19903 43821
rect 16589 43763 16594 43819
rect 16650 43763 19903 43819
rect 16589 43761 19903 43763
rect 16589 43758 16655 43761
rect 19903 43753 19967 43759
rect 17218 43669 17284 43672
rect 20099 43671 20163 43677
rect 17218 43667 20099 43669
rect 17218 43611 17223 43667
rect 17279 43611 20099 43667
rect 17218 43609 20099 43611
rect 17218 43606 17284 43609
rect 20099 43601 20163 43607
rect 18456 43526 18522 43529
rect 20621 43526 20627 43528
rect 18456 43524 20627 43526
rect 18456 43468 18461 43524
rect 18517 43468 20627 43524
rect 18456 43466 20627 43468
rect 18456 43463 18522 43466
rect 20621 43464 20627 43466
rect 20691 43464 20697 43528
rect 18166 43340 18232 43343
rect 20894 43342 20958 43348
rect 18166 43338 20894 43340
rect 18166 43282 18171 43338
rect 18227 43282 20894 43338
rect 18166 43280 20894 43282
rect 18166 43277 18232 43280
rect 9195 43271 9261 43276
rect 20894 43272 20958 43278
rect 9195 43215 9200 43271
rect 9256 43215 9261 43271
rect 9195 43210 9261 43215
rect 21650 43164 21716 43167
rect 25084 43166 25148 43172
rect 21650 43162 25084 43164
rect 20203 43150 20269 43153
rect 21408 43152 21472 43158
rect 20203 43148 21408 43150
rect 20203 43092 20208 43148
rect 20264 43092 21408 43148
rect 20203 43090 21408 43092
rect 20203 43087 20269 43090
rect 21650 43106 21655 43162
rect 21711 43106 25084 43162
rect 21650 43104 25084 43106
rect 21650 43101 21716 43104
rect 25084 43096 25148 43102
rect 21408 43082 21472 43088
rect 23553 42812 23619 42815
rect 25636 42814 25700 42820
rect 23553 42810 25636 42812
rect 23553 42754 23558 42810
rect 23614 42754 25636 42810
rect 23553 42752 25636 42754
rect 23553 42749 23619 42752
rect 25636 42744 25700 42750
rect 25948 32812 26008 44732
rect 23260 32752 26008 32812
rect 6160 21986 6560 24172
rect 192 21586 198 21986
rect 598 21586 26554 21986
rect 5630 21469 5842 21586
rect 5630 21267 5635 21469
rect 5837 21267 5842 21469
rect 5630 21262 5842 21267
rect 8430 21469 8642 21586
rect 8430 21267 8435 21469
rect 8637 21267 8642 21469
rect 8430 21262 8642 21267
rect 11230 21469 11442 21586
rect 11230 21267 11235 21469
rect 11437 21267 11442 21469
rect 11230 21262 11442 21267
rect 14030 21469 14242 21586
rect 14030 21267 14035 21469
rect 14237 21267 14242 21469
rect 14030 21262 14242 21267
rect 16830 21469 17042 21586
rect 16830 21267 16835 21469
rect 17037 21267 17042 21469
rect 19630 21469 19842 21586
rect 16830 21262 17042 21267
rect 17955 21364 18355 21370
rect 794 20634 800 21034
rect 1200 20964 17955 21034
rect 19630 21267 19635 21469
rect 19837 21267 19842 21469
rect 19630 21262 19842 21267
rect 22430 21469 22642 21586
rect 22430 21267 22435 21469
rect 22637 21267 22642 21469
rect 22430 21262 22642 21267
rect 25230 21469 25442 21586
rect 25230 21267 25235 21469
rect 25437 21267 25442 21469
rect 25230 21262 25442 21267
rect 18355 20964 26554 21034
rect 1200 20634 26554 20964
rect 4320 20527 4532 20634
rect 4320 20325 4325 20527
rect 4527 20325 4532 20527
rect 4320 20320 4532 20325
rect 7120 20527 7332 20634
rect 7120 20325 7125 20527
rect 7327 20325 7332 20527
rect 7120 20320 7332 20325
rect 9920 20527 10132 20634
rect 9920 20325 9925 20527
rect 10127 20325 10132 20527
rect 9920 20320 10132 20325
rect 12720 20527 12932 20634
rect 12720 20325 12725 20527
rect 12927 20325 12932 20527
rect 12720 20320 12932 20325
rect 15520 20527 15732 20634
rect 15520 20325 15525 20527
rect 15727 20325 15732 20527
rect 15520 20320 15732 20325
rect 18320 20527 18532 20634
rect 18320 20325 18325 20527
rect 18527 20325 18532 20527
rect 18320 20320 18532 20325
rect 21120 20527 21332 20634
rect 21120 20325 21125 20527
rect 21327 20325 21332 20527
rect 21120 20320 21332 20325
rect 23920 20527 24132 20634
rect 23920 20325 23925 20527
rect 24127 20325 24132 20527
rect 23920 20320 24132 20325
rect 6233 19763 6424 19764
rect 9033 19763 9224 19764
rect 11833 19763 12024 19764
rect 14633 19763 14824 19764
rect 17433 19763 17624 19764
rect 20233 19763 20424 19764
rect 23033 19763 23224 19764
rect 25833 19763 26024 19764
rect 6228 19574 6234 19763
rect 6423 19574 6429 19763
rect 9028 19574 9034 19763
rect 9223 19574 9229 19763
rect 11828 19574 11834 19763
rect 12023 19574 12029 19763
rect 14628 19574 14634 19763
rect 14823 19574 14829 19763
rect 17428 19574 17434 19763
rect 17623 19574 17629 19763
rect 20228 19574 20234 19763
rect 20423 19574 20429 19763
rect 23028 19574 23034 19763
rect 23223 19574 23229 19763
rect 25828 19574 25834 19763
rect 26023 19574 26029 19763
rect 6233 19521 6424 19574
rect 6233 19340 6238 19521
rect 6419 19340 6424 19521
rect 6233 19335 6424 19340
rect 9033 19521 9224 19574
rect 9033 19340 9038 19521
rect 9219 19340 9224 19521
rect 9033 19335 9224 19340
rect 11833 19521 12024 19574
rect 11833 19340 11838 19521
rect 12019 19340 12024 19521
rect 11833 19335 12024 19340
rect 14633 19521 14824 19574
rect 14633 19340 14638 19521
rect 14819 19340 14824 19521
rect 14633 19335 14824 19340
rect 17433 19521 17624 19574
rect 17433 19340 17438 19521
rect 17619 19340 17624 19521
rect 17433 19335 17624 19340
rect 20233 19521 20424 19574
rect 20233 19340 20238 19521
rect 20419 19340 20424 19521
rect 20233 19335 20424 19340
rect 23033 19521 23224 19574
rect 23033 19340 23038 19521
rect 23219 19340 23224 19521
rect 23033 19335 23224 19340
rect 25833 19521 26024 19574
rect 25833 19340 25838 19521
rect 26019 19340 26024 19521
rect 25833 19335 26024 19340
rect 801 2520 1199 2525
rect 800 2519 4964 2520
rect 800 2121 801 2519
rect 1199 2515 4964 2519
rect 1199 2125 4569 2515
rect 4959 2125 4964 2515
rect 1199 2121 4964 2125
rect 800 2120 4964 2121
rect 27169 2240 27474 2245
rect 801 2115 1199 2120
rect 27169 1945 27174 2240
rect 27469 1945 27474 2240
rect 27169 1940 27474 1945
rect 27174 1744 27469 1940
rect 27174 1443 27469 1449
<< via3 >>
rect 16654 44730 16718 44794
rect 8466 44568 8530 44632
rect 14189 44430 14253 44494
rect 14236 44282 14300 44346
rect 19514 44092 19578 44156
rect 19706 43916 19770 43980
rect 19903 43759 19967 43823
rect 20099 43607 20163 43671
rect 20627 43464 20691 43528
rect 20894 43278 20958 43342
rect 21408 43088 21472 43152
rect 25084 43102 25148 43166
rect 25636 42750 25700 42814
rect 198 21586 598 21986
rect 800 20634 1200 21034
rect 17955 20964 18355 21364
rect 6234 19574 6423 19763
rect 9034 19574 9223 19763
rect 11834 19574 12023 19763
rect 14634 19574 14823 19763
rect 17434 19574 17623 19763
rect 20234 19574 20423 19763
rect 23034 19574 23223 19763
rect 25834 19574 26023 19763
rect 801 2121 1199 2519
rect 27174 1449 27469 1744
<< metal4 >>
rect 3006 44792 3066 45152
rect 3558 44792 3618 45152
rect 4110 44792 4170 45152
rect 4662 44792 4722 45152
rect 5214 44792 5274 45152
rect 5766 44792 5826 45152
rect 6318 44792 6378 45152
rect 6870 44792 6930 45152
rect 7422 44792 7482 45152
rect 7974 44792 8034 45152
rect 8526 44792 8586 45152
rect 9078 44792 9138 45152
rect 9630 44792 9690 45152
rect 10182 44792 10242 45152
rect 10734 44792 10794 45152
rect 11286 44792 11346 45152
rect 11838 44792 11898 45152
rect 12390 44792 12450 45152
rect 12942 44792 13002 45152
rect 13494 44792 13554 45152
rect 14046 44792 14106 45152
rect 14598 44792 14658 45152
rect 15150 44792 15210 45152
rect 960 44732 15210 44792
rect 15702 44792 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44820 19626 45152
rect 16653 44794 16719 44795
rect 16653 44792 16654 44794
rect 15702 44732 16654 44792
rect 960 44152 1020 44732
rect 6870 44722 6930 44732
rect 7974 44716 8034 44732
rect 16653 44730 16654 44732
rect 16718 44730 16719 44794
rect 16653 44729 16719 44730
rect 18807 44760 19626 44820
rect 8465 44632 8531 44633
rect 8465 44568 8466 44632
rect 8530 44630 8531 44632
rect 18807 44630 18867 44760
rect 20118 44654 20178 45152
rect 8530 44570 18867 44630
rect 19103 44594 20178 44654
rect 8530 44568 8531 44570
rect 8465 44567 8531 44568
rect 14188 44494 14254 44495
rect 14188 44430 14189 44494
rect 14253 44492 14254 44494
rect 19103 44492 19163 44594
rect 20670 44501 20730 45152
rect 14253 44432 19163 44492
rect 19264 44441 20730 44501
rect 14253 44430 14254 44432
rect 14188 44429 14254 44430
rect 14235 44346 14301 44347
rect 14235 44282 14236 44346
rect 14300 44344 14301 44346
rect 19264 44344 19324 44441
rect 14300 44284 19324 44344
rect 21222 44325 21282 45152
rect 14300 44282 14301 44284
rect 14235 44281 14301 44282
rect 19516 44265 21282 44325
rect 19516 44157 19576 44265
rect 21774 44159 21834 45152
rect 19513 44156 19579 44157
rect 200 21987 600 44152
rect 197 21986 600 21987
rect 197 21586 198 21986
rect 598 21586 600 21986
rect 197 21585 600 21586
rect 200 1000 600 21585
rect 800 21035 1200 44152
rect 799 21034 1201 21035
rect 799 20634 800 21034
rect 1200 20634 1201 21034
rect 799 20633 1201 20634
rect 800 2519 1200 20633
rect 800 2121 801 2519
rect 1199 2121 1200 2519
rect 800 1000 1200 2121
rect 1400 20160 1800 44152
rect 19513 44092 19514 44156
rect 19578 44092 19579 44156
rect 19513 44091 19579 44092
rect 19708 44099 21834 44159
rect 19708 43981 19768 44099
rect 22326 44002 22386 45152
rect 19705 43980 19771 43981
rect 19705 43916 19706 43980
rect 19770 43916 19771 43980
rect 19705 43915 19771 43916
rect 19905 43942 22386 44002
rect 19905 43824 19965 43942
rect 22878 43845 22938 45152
rect 19902 43823 19968 43824
rect 19902 43759 19903 43823
rect 19967 43759 19968 43823
rect 19902 43758 19968 43759
rect 20101 43785 22938 43845
rect 20101 43672 20161 43785
rect 20098 43671 20164 43672
rect 20098 43607 20099 43671
rect 20163 43607 20164 43671
rect 23430 43669 23490 45152
rect 20098 43606 20164 43607
rect 20629 43609 23490 43669
rect 20629 43529 20689 43609
rect 20626 43528 20692 43529
rect 20626 43464 20627 43528
rect 20691 43464 20692 43528
rect 23982 43502 24042 45152
rect 20626 43463 20692 43464
rect 20896 43442 24042 43502
rect 20896 43343 20956 43442
rect 24534 43369 24594 45152
rect 20893 43342 20959 43343
rect 20893 43278 20894 43342
rect 20958 43278 20959 43342
rect 20893 43277 20959 43278
rect 21410 43309 24594 43369
rect 21410 43153 21470 43309
rect 25086 43167 25146 45152
rect 25083 43166 25149 43167
rect 21407 43152 21473 43153
rect 21407 43088 21408 43152
rect 21472 43088 21473 43152
rect 25083 43102 25084 43166
rect 25148 43102 25149 43166
rect 25083 43101 25149 43102
rect 21407 43087 21473 43088
rect 25638 42815 25698 45152
rect 26190 44952 26250 45152
rect 25635 42814 25701 42815
rect 25635 42750 25636 42814
rect 25700 42750 25701 42814
rect 25635 42749 25701 42750
rect 17955 21365 18355 24157
rect 17954 21364 18356 21365
rect 17954 20964 17955 21364
rect 18355 20964 18356 21364
rect 17954 20963 18356 20964
rect 1400 19763 26554 20160
rect 1400 19760 6234 19763
rect 1400 1000 1800 19760
rect 6233 19574 6234 19760
rect 6423 19760 9034 19763
rect 6423 19574 6424 19760
rect 6233 19573 6424 19574
rect 9033 19574 9034 19760
rect 9223 19760 11834 19763
rect 9223 19574 9224 19760
rect 9033 19573 9224 19574
rect 11833 19574 11834 19760
rect 12023 19760 14634 19763
rect 12023 19574 12024 19760
rect 11833 19573 12024 19574
rect 14633 19574 14634 19760
rect 14823 19760 17434 19763
rect 14823 19574 14824 19760
rect 14633 19573 14824 19574
rect 17433 19574 17434 19760
rect 17623 19760 20234 19763
rect 17623 19574 17624 19760
rect 17433 19573 17624 19574
rect 20233 19574 20234 19760
rect 20423 19760 23034 19763
rect 20423 19574 20424 19760
rect 20233 19573 20424 19574
rect 23033 19574 23034 19760
rect 23223 19760 25834 19763
rect 23223 19574 23224 19760
rect 23033 19573 23224 19574
rect 25833 19574 25834 19760
rect 26023 19760 26554 19763
rect 26023 19574 26024 19760
rect 25833 19573 26024 19574
rect 27173 1744 27470 1745
rect 27173 1449 27174 1744
rect 27469 1449 27470 1744
rect 27173 1448 27470 1449
rect 27174 315 27469 1448
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 0 27414 315
use dac_drive  dac_drive_1
array 0 0 -4800 0 7 2800
timestamp 1720097992
transform 0 1 5120 -1 0 16360
box -3000 -920 1360 1324
use r2r  r2r_0
timestamp 1720521779
transform 1 0 8664 0 -1 12768
box -1010 300 13300 11100
use r2r_dac_control  r2r_dac_control_0
timestamp 1720442423
transform 1 0 3433 0 1 22916
box 514 0 20000 20000
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1800 44152 1 FreeSans 1600 0 0 0 VAPWR
port 53 nsew power bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
