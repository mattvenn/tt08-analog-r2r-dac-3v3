magic
tech sky130A
magscale 1 2
timestamp 1720101481
<< viali >>
rect 3709 15045 3743 15079
rect 949 14977 983 15011
rect 1225 14977 1259 15011
rect 2237 14909 2271 14943
rect 3525 14909 3559 14943
rect 4537 14909 4571 14943
rect 4813 14909 4847 14943
rect 6101 14909 6135 14943
rect 7389 14909 7423 14943
rect 8677 14909 8711 14943
rect 9229 14909 9263 14943
rect 9965 14909 9999 14943
rect 11253 14909 11287 14943
rect 12541 14909 12575 14943
rect 13185 14909 13219 14943
rect 13921 14909 13955 14943
rect 2421 14773 2455 14807
rect 4629 14773 4663 14807
rect 4997 14773 5031 14807
rect 6285 14773 6319 14807
rect 7573 14773 7607 14807
rect 8861 14773 8895 14807
rect 9137 14773 9171 14807
rect 10149 14773 10183 14807
rect 11437 14773 11471 14807
rect 12725 14773 12759 14807
rect 13093 14773 13127 14807
rect 13645 14773 13679 14807
rect 14105 14773 14139 14807
rect 4629 14569 4663 14603
rect 9321 14569 9355 14603
rect 13185 14569 13219 14603
rect 13553 14501 13587 14535
rect 3516 14433 3550 14467
rect 5365 14433 5399 14467
rect 6009 14433 6043 14467
rect 6276 14433 6310 14467
rect 7481 14433 7515 14467
rect 7941 14433 7975 14467
rect 8208 14433 8242 14467
rect 9680 14433 9714 14467
rect 11621 14433 11655 14467
rect 11805 14433 11839 14467
rect 12061 14433 12095 14467
rect 3249 14365 3283 14399
rect 4721 14365 4755 14399
rect 5089 14365 5123 14399
rect 5181 14365 5215 14399
rect 9413 14365 9447 14399
rect 10977 14365 11011 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 13277 14365 13311 14399
rect 7389 14297 7423 14331
rect 7573 14229 7607 14263
rect 10793 14229 10827 14263
rect 15025 14229 15059 14263
rect 4537 14025 4571 14059
rect 4721 14025 4755 14059
rect 6285 14025 6319 14059
rect 6745 14025 6779 14059
rect 8033 14025 8067 14059
rect 9045 14025 9079 14059
rect 10425 14025 10459 14059
rect 10701 14025 10735 14059
rect 11897 14025 11931 14059
rect 12817 14025 12851 14059
rect 14197 14025 14231 14059
rect 5549 13957 5583 13991
rect 10885 13957 10919 13991
rect 6193 13889 6227 13923
rect 7941 13889 7975 13923
rect 8769 13889 8803 13923
rect 10425 13889 10459 13923
rect 4721 13821 4755 13855
rect 4905 13821 4939 13855
rect 5365 13821 5399 13855
rect 6101 13821 6135 13855
rect 6929 13821 6963 13855
rect 7021 13821 7055 13855
rect 7849 13821 7883 13855
rect 8861 13821 8895 13855
rect 10333 13821 10367 13855
rect 10793 13821 10827 13855
rect 11805 13821 11839 13855
rect 12081 13821 12115 13855
rect 12173 13821 12207 13855
rect 12817 13821 12851 13855
rect 13001 13821 13035 13855
rect 13277 13821 13311 13855
rect 13553 13821 13587 13855
rect 14105 13821 14139 13855
rect 6469 13685 6503 13719
rect 7389 13685 7423 13719
rect 8217 13685 8251 13719
rect 8401 13685 8435 13719
rect 11621 13685 11655 13719
rect 12541 13685 12575 13719
rect 12633 13685 12667 13719
rect 13093 13685 13127 13719
rect 13645 13685 13679 13719
rect 5089 13481 5123 13515
rect 5181 13481 5215 13515
rect 7389 13481 7423 13515
rect 6070 13413 6104 13447
rect 10701 13413 10735 13447
rect 15025 13413 15059 13447
rect 3821 13345 3855 13379
rect 4077 13345 4111 13379
rect 4721 13345 4755 13379
rect 5365 13345 5399 13379
rect 5549 13345 5583 13379
rect 5825 13345 5859 13379
rect 7665 13345 7699 13379
rect 7757 13345 7791 13379
rect 8677 13345 8711 13379
rect 9404 13345 9438 13379
rect 10609 13345 10643 13379
rect 11529 13345 11563 13379
rect 13001 13345 13035 13379
rect 13645 13345 13679 13379
rect 4445 13277 4479 13311
rect 4629 13277 4663 13311
rect 8769 13277 8803 13311
rect 9137 13277 9171 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 10517 13209 10551 13243
rect 2697 13141 2731 13175
rect 5365 13141 5399 13175
rect 7205 13141 7239 13175
rect 7573 13141 7607 13175
rect 8861 13141 8895 13175
rect 9045 13141 9079 13175
rect 11437 13141 11471 13175
rect 11897 13141 11931 13175
rect 4905 12937 4939 12971
rect 5825 12937 5859 12971
rect 6837 12937 6871 12971
rect 9873 12937 9907 12971
rect 11897 12937 11931 12971
rect 8677 12869 8711 12903
rect 6101 12801 6135 12835
rect 6469 12801 6503 12835
rect 9229 12801 9263 12835
rect 9597 12801 9631 12835
rect 11529 12801 11563 12835
rect 12081 12801 12115 12835
rect 12449 12801 12483 12835
rect 12817 12801 12851 12835
rect 13829 12801 13863 12835
rect 4169 12733 4203 12767
rect 4353 12733 4387 12767
rect 4537 12733 4571 12767
rect 4813 12733 4847 12767
rect 6009 12733 6043 12767
rect 6929 12733 6963 12767
rect 9689 12733 9723 12767
rect 11713 12733 11747 12767
rect 12357 12733 12391 12767
rect 13001 12733 13035 12767
rect 13185 12733 13219 12767
rect 13921 12733 13955 12767
rect 4445 12665 4479 12699
rect 8401 12665 8435 12699
rect 11989 12665 12023 12699
rect 4721 12597 4755 12631
rect 8861 12597 8895 12631
rect 12633 12597 12667 12631
rect 13553 12597 13587 12631
rect 4629 12393 4663 12427
rect 11345 12393 11379 12427
rect 11713 12393 11747 12427
rect 4261 12325 4295 12359
rect 4721 12325 4755 12359
rect 7113 12325 7147 12359
rect 7481 12325 7515 12359
rect 11253 12325 11287 12359
rect 3617 12257 3651 12291
rect 3985 12257 4019 12291
rect 4133 12257 4167 12291
rect 4353 12257 4387 12291
rect 4450 12257 4484 12291
rect 4905 12257 4939 12291
rect 5181 12257 5215 12291
rect 5365 12257 5399 12291
rect 6837 12257 6871 12291
rect 7021 12257 7055 12291
rect 7205 12257 7239 12291
rect 7665 12257 7699 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8309 12257 8343 12291
rect 8401 12257 8435 12291
rect 8585 12257 8619 12291
rect 8677 12257 8711 12291
rect 8769 12257 8803 12291
rect 11805 12257 11839 12291
rect 7849 12189 7883 12223
rect 7941 12189 7975 12223
rect 11161 12189 11195 12223
rect 7389 12121 7423 12155
rect 8953 12121 8987 12155
rect 3801 12053 3835 12087
rect 13093 12053 13127 12087
rect 4353 11849 4387 11883
rect 7389 11849 7423 11883
rect 8493 11849 8527 11883
rect 12633 11849 12667 11883
rect 12725 11849 12759 11883
rect 4813 11781 4847 11815
rect 5181 11781 5215 11815
rect 4905 11713 4939 11747
rect 10333 11713 10367 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 12541 11713 12575 11747
rect 4261 11645 4295 11679
rect 4537 11645 4571 11679
rect 4629 11645 4663 11679
rect 8769 11645 8803 11679
rect 8861 11645 8895 11679
rect 8953 11645 8987 11679
rect 9137 11645 9171 11679
rect 9597 11645 9631 11679
rect 9781 11645 9815 11679
rect 9873 11645 9907 11679
rect 9965 11645 9999 11679
rect 10149 11645 10183 11679
rect 10793 11645 10827 11679
rect 11345 11645 11379 11679
rect 11713 11645 11747 11679
rect 12173 11645 12207 11679
rect 12817 11645 12851 11679
rect 13553 11645 13587 11679
rect 13737 11645 13771 11679
rect 6101 11577 6135 11611
rect 5365 11509 5399 11543
rect 10425 11509 10459 11543
rect 11529 11509 11563 11543
rect 11805 11509 11839 11543
rect 12265 11509 12299 11543
rect 13645 11509 13679 11543
rect 7757 11305 7791 11339
rect 8493 11305 8527 11339
rect 9597 11305 9631 11339
rect 11713 11305 11747 11339
rect 13277 11305 13311 11339
rect 6092 11237 6126 11271
rect 8861 11237 8895 11271
rect 10425 11237 10459 11271
rect 5181 11169 5215 11203
rect 5365 11169 5399 11203
rect 5825 11169 5859 11203
rect 7297 11169 7331 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 8677 11169 8711 11203
rect 8769 11169 8803 11203
rect 9045 11169 9079 11203
rect 9781 11169 9815 11203
rect 9873 11169 9907 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 10977 11169 11011 11203
rect 11161 11169 11195 11203
rect 11805 11169 11839 11203
rect 12541 11169 12575 11203
rect 12725 11169 12759 11203
rect 12817 11169 12851 11203
rect 13093 11169 13127 11203
rect 11621 11101 11655 11135
rect 12909 11101 12943 11135
rect 13369 11101 13403 11135
rect 13645 11101 13679 11135
rect 5365 10965 5399 10999
rect 7205 10965 7239 10999
rect 7389 10965 7423 10999
rect 7941 10965 7975 10999
rect 10333 10965 10367 10999
rect 11069 10965 11103 10999
rect 12173 10965 12207 10999
rect 14933 10965 14967 10999
rect 6193 10761 6227 10795
rect 6469 10761 6503 10795
rect 12817 10761 12851 10795
rect 13001 10761 13035 10795
rect 6561 10693 6595 10727
rect 9689 10693 9723 10727
rect 14289 10693 14323 10727
rect 4629 10625 4663 10659
rect 5365 10625 5399 10659
rect 5733 10625 5767 10659
rect 6653 10625 6687 10659
rect 9321 10625 9355 10659
rect 11621 10625 11655 10659
rect 11989 10625 12023 10659
rect 14933 10625 14967 10659
rect 5457 10557 5491 10591
rect 5641 10557 5675 10591
rect 5825 10557 5859 10591
rect 6009 10557 6043 10591
rect 6377 10557 6411 10591
rect 9137 10557 9171 10591
rect 9413 10557 9447 10591
rect 11529 10557 11563 10591
rect 12081 10557 12115 10591
rect 12265 10557 12299 10591
rect 12541 10557 12575 10591
rect 13553 10557 13587 10591
rect 14197 10557 14231 10591
rect 4384 10489 4418 10523
rect 9505 10489 9539 10523
rect 9689 10489 9723 10523
rect 11345 10489 11379 10523
rect 13185 10489 13219 10523
rect 3249 10421 3283 10455
rect 4721 10421 4755 10455
rect 8953 10421 8987 10455
rect 11713 10421 11747 10455
rect 11897 10421 11931 10455
rect 12725 10421 12759 10455
rect 12985 10421 13019 10455
rect 4721 10217 4755 10251
rect 5825 10217 5859 10251
rect 6193 10217 6227 10251
rect 7021 10217 7055 10251
rect 8493 10217 8527 10251
rect 10609 10217 10643 10251
rect 6377 10149 6411 10183
rect 7358 10149 7392 10183
rect 11253 10149 11287 10183
rect 11805 10149 11839 10183
rect 12021 10149 12055 10183
rect 12265 10149 12299 10183
rect 12449 10149 12483 10183
rect 12633 10149 12667 10183
rect 14657 10149 14691 10183
rect 4445 10081 4479 10115
rect 4905 10081 4939 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 6009 10081 6043 10115
rect 6101 10081 6135 10115
rect 6837 10081 6871 10115
rect 8769 10081 8803 10115
rect 8953 10081 8987 10115
rect 9045 10081 9079 10115
rect 9229 10081 9263 10115
rect 9496 10081 9530 10115
rect 11437 10081 11471 10115
rect 11621 10081 11655 10115
rect 13001 10081 13035 10115
rect 4261 10013 4295 10047
rect 4629 10013 4663 10047
rect 5089 10013 5123 10047
rect 5181 10013 5215 10047
rect 7113 10013 7147 10047
rect 11713 10013 11747 10047
rect 13277 10013 13311 10047
rect 12173 9945 12207 9979
rect 8585 9877 8619 9911
rect 11529 9877 11563 9911
rect 11989 9877 12023 9911
rect 5089 9673 5123 9707
rect 6285 9673 6319 9707
rect 11621 9673 11655 9707
rect 6101 9605 6135 9639
rect 8217 9605 8251 9639
rect 6009 9537 6043 9571
rect 7389 9537 7423 9571
rect 9229 9537 9263 9571
rect 5549 9469 5583 9503
rect 5641 9469 5675 9503
rect 7021 9469 7055 9503
rect 7113 9469 7147 9503
rect 7481 9469 7515 9503
rect 8033 9469 8067 9503
rect 10977 9469 11011 9503
rect 11345 9469 11379 9503
rect 11621 9469 11655 9503
rect 12817 9469 12851 9503
rect 13001 9469 13035 9503
rect 13553 9469 13587 9503
rect 13737 9469 13771 9503
rect 13921 9469 13955 9503
rect 5273 9401 5307 9435
rect 5917 9401 5951 9435
rect 6469 9401 6503 9435
rect 7849 9401 7883 9435
rect 4905 9333 4939 9367
rect 5073 9333 5107 9367
rect 5365 9333 5399 9367
rect 6269 9333 6303 9367
rect 6837 9333 6871 9367
rect 7665 9333 7699 9367
rect 7941 9333 7975 9367
rect 11437 9333 11471 9367
rect 12633 9333 12667 9367
rect 4721 9129 4755 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 7087 9129 7121 9163
rect 9689 9129 9723 9163
rect 10701 9129 10735 9163
rect 7297 9061 7331 9095
rect 11805 9061 11839 9095
rect 13277 9061 13311 9095
rect 3608 8993 3642 9027
rect 5273 8993 5307 9027
rect 5549 8993 5583 9027
rect 8953 8993 8987 9027
rect 9137 8993 9171 9027
rect 9229 8993 9263 9027
rect 9321 8993 9355 9027
rect 9505 8993 9539 9027
rect 10517 8993 10551 9027
rect 11345 8993 11379 9027
rect 11437 8993 11471 9027
rect 12541 8993 12575 9027
rect 12725 8993 12759 9027
rect 13093 8993 13127 9027
rect 13645 8993 13679 9027
rect 3341 8925 3375 8959
rect 10977 8925 11011 8959
rect 11621 8925 11655 8959
rect 12817 8925 12851 8959
rect 12909 8925 12943 8959
rect 13369 8925 13403 8959
rect 6929 8857 6963 8891
rect 7113 8789 7147 8823
rect 11897 8789 11931 8823
rect 14933 8789 14967 8823
rect 3709 8585 3743 8619
rect 5365 8585 5399 8619
rect 6929 8585 6963 8619
rect 9137 8585 9171 8619
rect 13553 8585 13587 8619
rect 11437 8517 11471 8551
rect 11713 8517 11747 8551
rect 11897 8517 11931 8551
rect 8401 8449 8435 8483
rect 8493 8449 8527 8483
rect 11529 8449 11563 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 3893 8381 3927 8415
rect 3985 8381 4019 8415
rect 6469 8381 6503 8415
rect 6561 8381 6595 8415
rect 6653 8381 6687 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 7297 8381 7331 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 8769 8381 8803 8415
rect 8861 8381 8895 8415
rect 10517 8381 10551 8415
rect 11161 8381 11195 8415
rect 11805 8381 11839 8415
rect 13737 8381 13771 8415
rect 14013 8381 14047 8415
rect 14197 8381 14231 8415
rect 4252 8313 4286 8347
rect 6193 8313 6227 8347
rect 7849 8313 7883 8347
rect 10250 8313 10284 8347
rect 11437 8313 11471 8347
rect 11529 8313 11563 8347
rect 8217 8245 8251 8279
rect 9045 8245 9079 8279
rect 11253 8245 11287 8279
rect 12265 8245 12299 8279
rect 7915 8041 7949 8075
rect 8509 8041 8543 8075
rect 8677 8041 8711 8075
rect 9413 8041 9447 8075
rect 7665 7973 7699 8007
rect 8125 7973 8159 8007
rect 8309 7973 8343 8007
rect 8795 7973 8829 8007
rect 8985 7973 9019 8007
rect 9229 7905 9263 7939
rect 10425 7905 10459 7939
rect 13645 7905 13679 7939
rect 13369 7837 13403 7871
rect 9137 7769 9171 7803
rect 6193 7701 6227 7735
rect 7757 7701 7791 7735
rect 7941 7701 7975 7735
rect 8493 7701 8527 7735
rect 8953 7701 8987 7735
rect 10517 7701 10551 7735
rect 14749 7701 14783 7735
rect 5825 7497 5859 7531
rect 6561 7497 6595 7531
rect 7757 7429 7791 7463
rect 12909 7429 12943 7463
rect 6745 7361 6779 7395
rect 7113 7361 7147 7395
rect 7205 7361 7239 7395
rect 14105 7361 14139 7395
rect 5641 7293 5675 7327
rect 6377 7293 6411 7327
rect 6837 7293 6871 7327
rect 7941 7293 7975 7327
rect 8033 7293 8067 7327
rect 11345 7293 11379 7327
rect 11529 7293 11563 7327
rect 11621 7293 11655 7327
rect 13921 7293 13955 7327
rect 6009 7225 6043 7259
rect 6101 7225 6135 7259
rect 7757 7225 7791 7259
rect 5089 7157 5123 7191
rect 6193 7157 6227 7191
rect 11529 7157 11563 7191
rect 13553 7157 13587 7191
rect 14013 7157 14047 7191
rect 5825 6953 5859 6987
rect 6761 6953 6795 6987
rect 6929 6953 6963 6987
rect 9781 6953 9815 6987
rect 10977 6953 11011 6987
rect 11437 6953 11471 6987
rect 6377 6885 6411 6919
rect 6561 6885 6595 6919
rect 8309 6885 8343 6919
rect 8646 6885 8680 6919
rect 13553 6885 13587 6919
rect 3700 6817 3734 6851
rect 5273 6817 5307 6851
rect 5365 6817 5399 6851
rect 5457 6820 5491 6854
rect 5641 6817 5675 6851
rect 6009 6817 6043 6851
rect 6101 6817 6135 6851
rect 7573 6817 7607 6851
rect 7757 6817 7791 6851
rect 7941 6817 7975 6851
rect 8125 6817 8159 6851
rect 10149 6817 10183 6851
rect 10333 6817 10367 6851
rect 11345 6817 11379 6851
rect 12173 6817 12207 6851
rect 12541 6817 12575 6851
rect 12725 6817 12759 6851
rect 12909 6817 12943 6851
rect 13001 6817 13035 6851
rect 13461 6817 13495 6851
rect 3433 6749 3467 6783
rect 4997 6749 5031 6783
rect 6469 6749 6503 6783
rect 7849 6749 7883 6783
rect 8401 6749 8435 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 12081 6749 12115 6783
rect 12265 6749 12299 6783
rect 13185 6749 13219 6783
rect 13277 6681 13311 6715
rect 4813 6613 4847 6647
rect 6745 6613 6779 6647
rect 10333 6613 10367 6647
rect 12449 6613 12483 6647
rect 13093 6613 13127 6647
rect 7297 6409 7331 6443
rect 7665 6409 7699 6443
rect 12725 6409 12759 6443
rect 13185 6409 13219 6443
rect 13369 6409 13403 6443
rect 4813 6341 4847 6375
rect 5641 6273 5675 6307
rect 6561 6273 6595 6307
rect 8033 6273 8067 6307
rect 3433 6205 3467 6239
rect 5733 6205 5767 6239
rect 6193 6205 6227 6239
rect 6377 6205 6411 6239
rect 7113 6205 7147 6239
rect 7849 6205 7883 6239
rect 9781 6205 9815 6239
rect 12449 6205 12483 6239
rect 12725 6205 12759 6239
rect 13829 6205 13863 6239
rect 14473 6205 14507 6239
rect 3700 6137 3734 6171
rect 6009 6137 6043 6171
rect 6101 6137 6135 6171
rect 10048 6137 10082 6171
rect 13001 6137 13035 6171
rect 5457 6069 5491 6103
rect 11161 6069 11195 6103
rect 12541 6069 12575 6103
rect 13201 6069 13235 6103
rect 9597 5865 9631 5899
rect 11897 5865 11931 5899
rect 7573 5797 7607 5831
rect 8661 5797 8695 5831
rect 8861 5797 8895 5831
rect 9873 5797 9907 5831
rect 5641 5729 5675 5763
rect 6377 5729 6411 5763
rect 6469 5729 6503 5763
rect 7757 5729 7791 5763
rect 7849 5729 7883 5763
rect 8033 5729 8067 5763
rect 9781 5729 9815 5763
rect 9965 5729 9999 5763
rect 11713 5729 11747 5763
rect 12725 5729 12759 5763
rect 13001 5729 13035 5763
rect 13185 5729 13219 5763
rect 13369 5729 13403 5763
rect 13645 5661 13679 5695
rect 8493 5593 8527 5627
rect 10149 5593 10183 5627
rect 4997 5525 5031 5559
rect 6653 5525 6687 5559
rect 7573 5525 7607 5559
rect 8217 5525 8251 5559
rect 8677 5525 8711 5559
rect 12541 5525 12575 5559
rect 14933 5525 14967 5559
rect 4905 5321 4939 5355
rect 10057 5321 10091 5355
rect 12817 5321 12851 5355
rect 13185 5321 13219 5355
rect 9781 5253 9815 5287
rect 10241 5253 10275 5287
rect 12541 5253 12575 5287
rect 6285 5185 6319 5219
rect 7021 5185 7055 5219
rect 8125 5185 8159 5219
rect 8401 5185 8435 5219
rect 10977 5185 11011 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12725 5185 12759 5219
rect 14013 5185 14047 5219
rect 14565 5185 14599 5219
rect 5181 5117 5215 5151
rect 5273 5117 5307 5151
rect 5365 5117 5399 5151
rect 5549 5117 5583 5151
rect 5825 5117 5859 5151
rect 5917 5117 5951 5151
rect 6745 5117 6779 5151
rect 6929 5117 6963 5151
rect 7159 5117 7193 5151
rect 7297 5117 7331 5151
rect 7573 5117 7607 5151
rect 8657 5117 8691 5151
rect 10517 5117 10551 5151
rect 10609 5117 10643 5151
rect 11437 5117 11471 5151
rect 11621 5117 11655 5151
rect 12000 5117 12034 5151
rect 12265 5117 12299 5151
rect 13001 5117 13035 5151
rect 6193 5049 6227 5083
rect 9873 5049 9907 5083
rect 10089 5049 10123 5083
rect 10885 5049 10919 5083
rect 12357 5049 12391 5083
rect 12541 5049 12575 5083
rect 5641 4981 5675 5015
rect 7481 4981 7515 5015
rect 10333 4981 10367 5015
rect 12173 4981 12207 5015
rect 5457 4777 5491 4811
rect 6193 4777 6227 4811
rect 6745 4777 6779 4811
rect 8677 4777 8711 4811
rect 9413 4777 9447 4811
rect 10609 4777 10643 4811
rect 11713 4777 11747 4811
rect 14657 4777 14691 4811
rect 7858 4709 7892 4743
rect 12918 4709 12952 4743
rect 4077 4641 4111 4675
rect 4344 4641 4378 4675
rect 6009 4641 6043 4675
rect 6285 4641 6319 4675
rect 8125 4641 8159 4675
rect 8953 4641 8987 4675
rect 9321 4641 9355 4675
rect 9597 4641 9631 4675
rect 10425 4641 10459 4675
rect 10701 4641 10735 4675
rect 11345 4641 11379 4675
rect 11529 4641 11563 4675
rect 13185 4641 13219 4675
rect 13277 4641 13311 4675
rect 13553 4641 13587 4675
rect 8861 4573 8895 4607
rect 9229 4573 9263 4607
rect 9689 4573 9723 4607
rect 9781 4573 9815 4607
rect 9873 4573 9907 4607
rect 11805 4505 11839 4539
rect 5825 4437 5859 4471
rect 10241 4437 10275 4471
rect 4445 4233 4479 4267
rect 5181 4233 5215 4267
rect 6101 4233 6135 4267
rect 10241 4233 10275 4267
rect 4629 4029 4663 4063
rect 5365 3961 5399 3995
rect 5917 3961 5951 3995
rect 6133 3961 6167 3995
rect 10057 3961 10091 3995
rect 10273 3961 10307 3995
rect 4997 3893 5031 3927
rect 5165 3893 5199 3927
rect 6285 3893 6319 3927
rect 10425 3893 10459 3927
rect 10793 3689 10827 3723
rect 9413 3553 9447 3587
rect 9680 3553 9714 3587
rect 10057 3145 10091 3179
rect 10241 2941 10275 2975
<< metal1 >>
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 3697 15079 3755 15085
rect 3697 15045 3709 15079
rect 3743 15076 3755 15079
rect 5074 15076 5080 15088
rect 3743 15048 5080 15076
rect 3743 15045 3755 15048
rect 3697 15039 3755 15045
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 934 14968 940 15020
rect 992 14968 998 15020
rect 1213 15011 1271 15017
rect 1213 14977 1225 15011
rect 1259 15008 1271 15011
rect 4430 15008 4436 15020
rect 1259 14980 4436 15008
rect 1259 14977 1271 14980
rect 1213 14971 1271 14977
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 2130 14900 2136 14952
rect 2188 14940 2194 14952
rect 2225 14943 2283 14949
rect 2225 14940 2237 14943
rect 2188 14912 2237 14940
rect 2188 14900 2194 14912
rect 2225 14909 2237 14912
rect 2271 14909 2283 14943
rect 2225 14903 2283 14909
rect 3510 14900 3516 14952
rect 3568 14900 3574 14952
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4614 14940 4620 14952
rect 4571 14912 4620 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 4798 14900 4804 14952
rect 4856 14900 4862 14952
rect 5810 14900 5816 14952
rect 5868 14940 5874 14952
rect 6089 14943 6147 14949
rect 6089 14940 6101 14943
rect 5868 14912 6101 14940
rect 5868 14900 5874 14912
rect 6089 14909 6101 14912
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 7282 14900 7288 14952
rect 7340 14940 7346 14952
rect 7377 14943 7435 14949
rect 7377 14940 7389 14943
rect 7340 14912 7389 14940
rect 7340 14900 7346 14912
rect 7377 14909 7389 14912
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 9214 14900 9220 14952
rect 9272 14900 9278 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14940 10011 14943
rect 10042 14940 10048 14952
rect 9999 14912 10048 14940
rect 9999 14909 10011 14912
rect 9953 14903 10011 14909
rect 10042 14900 10048 14912
rect 10100 14900 10106 14952
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 11204 14912 11253 14940
rect 11204 14900 11210 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12529 14943 12587 14949
rect 12529 14940 12541 14943
rect 12492 14912 12541 14940
rect 12492 14900 12498 14912
rect 12529 14909 12541 14912
rect 12575 14909 12587 14943
rect 12529 14903 12587 14909
rect 13170 14900 13176 14952
rect 13228 14900 13234 14952
rect 13722 14900 13728 14952
rect 13780 14940 13786 14952
rect 13909 14943 13967 14949
rect 13909 14940 13921 14943
rect 13780 14912 13921 14940
rect 13780 14900 13786 14912
rect 13909 14909 13921 14912
rect 13955 14909 13967 14943
rect 13909 14903 13967 14909
rect 2409 14807 2467 14813
rect 2409 14773 2421 14807
rect 2455 14804 2467 14807
rect 3602 14804 3608 14816
rect 2455 14776 3608 14804
rect 2455 14773 2467 14776
rect 2409 14767 2467 14773
rect 3602 14764 3608 14776
rect 3660 14764 3666 14816
rect 4617 14807 4675 14813
rect 4617 14773 4629 14807
rect 4663 14804 4675 14807
rect 4706 14804 4712 14816
rect 4663 14776 4712 14804
rect 4663 14773 4675 14776
rect 4617 14767 4675 14773
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 4982 14764 4988 14816
rect 5040 14764 5046 14816
rect 6273 14807 6331 14813
rect 6273 14773 6285 14807
rect 6319 14804 6331 14807
rect 6362 14804 6368 14816
rect 6319 14776 6368 14804
rect 6319 14773 6331 14776
rect 6273 14767 6331 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 6972 14776 7573 14804
rect 6972 14764 6978 14776
rect 7561 14773 7573 14776
rect 7607 14773 7619 14807
rect 7561 14767 7619 14773
rect 8846 14764 8852 14816
rect 8904 14764 8910 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8996 14776 9137 14804
rect 8996 14764 9002 14776
rect 9125 14773 9137 14776
rect 9171 14773 9183 14807
rect 9125 14767 9183 14773
rect 10137 14807 10195 14813
rect 10137 14773 10149 14807
rect 10183 14804 10195 14807
rect 10410 14804 10416 14816
rect 10183 14776 10416 14804
rect 10183 14773 10195 14776
rect 10137 14767 10195 14773
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 11422 14764 11428 14816
rect 11480 14764 11486 14816
rect 12710 14764 12716 14816
rect 12768 14764 12774 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13081 14807 13139 14813
rect 13081 14804 13093 14807
rect 12860 14776 13093 14804
rect 12860 14764 12866 14776
rect 13081 14773 13093 14776
rect 13127 14773 13139 14807
rect 13081 14767 13139 14773
rect 13630 14764 13636 14816
rect 13688 14764 13694 14816
rect 14090 14764 14096 14816
rect 14148 14764 14154 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 4614 14560 4620 14612
rect 4672 14560 4678 14612
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9309 14603 9367 14609
rect 9309 14600 9321 14603
rect 9272 14572 9321 14600
rect 9272 14560 9278 14572
rect 9309 14569 9321 14572
rect 9355 14569 9367 14603
rect 9309 14563 9367 14569
rect 13170 14560 13176 14612
rect 13228 14560 13234 14612
rect 7374 14532 7380 14544
rect 6012 14504 7380 14532
rect 3504 14467 3562 14473
rect 3504 14433 3516 14467
rect 3550 14464 3562 14467
rect 5353 14467 5411 14473
rect 5353 14464 5365 14467
rect 3550 14436 5365 14464
rect 3550 14433 3562 14436
rect 3504 14427 3562 14433
rect 5353 14433 5365 14436
rect 5399 14433 5411 14467
rect 5810 14464 5816 14476
rect 5353 14427 5411 14433
rect 5506 14436 5816 14464
rect 3234 14356 3240 14408
rect 3292 14356 3298 14408
rect 4522 14356 4528 14408
rect 4580 14396 4586 14408
rect 4709 14399 4767 14405
rect 4709 14396 4721 14399
rect 4580 14368 4721 14396
rect 4580 14356 4586 14368
rect 4709 14365 4721 14368
rect 4755 14365 4767 14399
rect 4709 14359 4767 14365
rect 5074 14356 5080 14408
rect 5132 14356 5138 14408
rect 5166 14356 5172 14408
rect 5224 14356 5230 14408
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 5506 14260 5534 14436
rect 5810 14424 5816 14436
rect 5868 14464 5874 14476
rect 6012 14473 6040 14504
rect 7374 14492 7380 14504
rect 7432 14532 7438 14544
rect 13541 14535 13599 14541
rect 7432 14504 7972 14532
rect 7432 14492 7438 14504
rect 5997 14467 6055 14473
rect 5997 14464 6009 14467
rect 5868 14436 6009 14464
rect 5868 14424 5874 14436
rect 5997 14433 6009 14436
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6264 14467 6322 14473
rect 6264 14433 6276 14467
rect 6310 14464 6322 14467
rect 6730 14464 6736 14476
rect 6310 14436 6736 14464
rect 6310 14433 6322 14436
rect 6264 14427 6322 14433
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 7944 14473 7972 14504
rect 9416 14504 11836 14532
rect 7469 14467 7527 14473
rect 7469 14464 7481 14467
rect 7392 14436 7481 14464
rect 7392 14337 7420 14436
rect 7469 14433 7481 14436
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 7929 14467 7987 14473
rect 7929 14433 7941 14467
rect 7975 14433 7987 14467
rect 7929 14427 7987 14433
rect 8196 14467 8254 14473
rect 8196 14433 8208 14467
rect 8242 14464 8254 14467
rect 9030 14464 9036 14476
rect 8242 14436 9036 14464
rect 8242 14433 8254 14436
rect 8196 14427 8254 14433
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9416 14405 9444 14504
rect 11808 14473 11836 14504
rect 13541 14501 13553 14535
rect 13587 14532 13599 14535
rect 13630 14532 13636 14544
rect 13587 14504 13636 14532
rect 13587 14501 13599 14504
rect 13541 14495 13599 14501
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 14182 14492 14188 14544
rect 14240 14492 14246 14544
rect 9668 14467 9726 14473
rect 9668 14433 9680 14467
rect 9714 14464 9726 14467
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 9714 14436 11621 14464
rect 9714 14433 9726 14436
rect 9668 14427 9726 14433
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 11609 14427 11667 14433
rect 11793 14467 11851 14473
rect 11793 14433 11805 14467
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 12049 14467 12107 14473
rect 12049 14464 12061 14467
rect 11940 14436 12061 14464
rect 11940 14424 11946 14436
rect 12049 14433 12061 14436
rect 12095 14433 12107 14467
rect 12049 14427 12107 14433
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9180 14368 9413 14396
rect 9180 14356 9186 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11238 14356 11244 14408
rect 11296 14396 11302 14408
rect 11333 14399 11391 14405
rect 11333 14396 11345 14399
rect 11296 14368 11345 14396
rect 11296 14356 11302 14368
rect 11333 14365 11345 14368
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13136 14368 13277 14396
rect 13136 14356 13142 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 7377 14331 7435 14337
rect 7377 14297 7389 14331
rect 7423 14297 7435 14331
rect 7377 14291 7435 14297
rect 3292 14232 5534 14260
rect 3292 14220 3298 14232
rect 7558 14220 7564 14272
rect 7616 14220 7622 14272
rect 10778 14220 10784 14272
rect 10836 14220 10842 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 15013 14263 15071 14269
rect 15013 14260 15025 14263
rect 11848 14232 15025 14260
rect 11848 14220 11854 14232
rect 15013 14229 15025 14232
rect 15059 14229 15071 14263
rect 15013 14223 15071 14229
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 4522 14016 4528 14068
rect 4580 14016 4586 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 6270 14016 6276 14068
rect 6328 14016 6334 14068
rect 6730 14016 6736 14068
rect 6788 14016 6794 14068
rect 8021 14059 8079 14065
rect 8021 14025 8033 14059
rect 8067 14056 8079 14059
rect 8386 14056 8392 14068
rect 8067 14028 8392 14056
rect 8067 14025 8079 14028
rect 8021 14019 8079 14025
rect 8386 14016 8392 14028
rect 8444 14056 8450 14068
rect 8938 14056 8944 14068
rect 8444 14028 8944 14056
rect 8444 14016 8450 14028
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 9030 14016 9036 14068
rect 9088 14016 9094 14068
rect 10413 14059 10471 14065
rect 10413 14025 10425 14059
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 10689 14059 10747 14065
rect 10689 14025 10701 14059
rect 10735 14056 10747 14059
rect 10962 14056 10968 14068
rect 10735 14028 10968 14056
rect 10735 14025 10747 14028
rect 10689 14019 10747 14025
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 5224 13960 5549 13988
rect 5224 13948 5230 13960
rect 5537 13957 5549 13960
rect 5583 13988 5595 13991
rect 7006 13988 7012 14000
rect 5583 13960 7012 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 7006 13948 7012 13960
rect 7064 13988 7070 14000
rect 10428 13988 10456 14019
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11882 14016 11888 14068
rect 11940 14016 11946 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12802 14056 12808 14068
rect 12032 14028 12808 14056
rect 12032 14016 12038 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 14182 14016 14188 14068
rect 14240 14016 14246 14068
rect 10502 13988 10508 14000
rect 7064 13960 8800 13988
rect 10428 13960 10508 13988
rect 7064 13948 7070 13960
rect 5626 13920 5632 13932
rect 4908 13892 5632 13920
rect 4430 13812 4436 13864
rect 4488 13852 4494 13864
rect 4908 13861 4936 13892
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 6181 13923 6239 13929
rect 6181 13920 6193 13923
rect 6012 13892 6193 13920
rect 4709 13855 4767 13861
rect 4709 13852 4721 13855
rect 4488 13824 4721 13852
rect 4488 13812 4494 13824
rect 4709 13821 4721 13824
rect 4755 13821 4767 13855
rect 4709 13815 4767 13821
rect 4893 13855 4951 13861
rect 4893 13821 4905 13855
rect 4939 13821 4951 13855
rect 5353 13855 5411 13861
rect 5353 13852 5365 13855
rect 4893 13815 4951 13821
rect 5276 13824 5365 13852
rect 4724 13784 4752 13815
rect 5276 13796 5304 13824
rect 5353 13821 5365 13824
rect 5399 13852 5411 13855
rect 6012 13852 6040 13892
rect 6181 13889 6193 13892
rect 6227 13920 6239 13923
rect 7650 13920 7656 13932
rect 6227 13892 7656 13920
rect 6227 13889 6239 13892
rect 6181 13883 6239 13889
rect 7650 13880 7656 13892
rect 7708 13920 7714 13932
rect 8772 13929 8800 13960
rect 10502 13948 10508 13960
rect 10560 13988 10566 14000
rect 10873 13991 10931 13997
rect 10873 13988 10885 13991
rect 10560 13960 10885 13988
rect 10560 13948 10566 13960
rect 10873 13957 10885 13960
rect 10919 13957 10931 13991
rect 10873 13951 10931 13957
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7708 13892 7941 13920
rect 7708 13880 7714 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8757 13923 8815 13929
rect 8757 13889 8769 13923
rect 8803 13920 8815 13923
rect 9490 13920 9496 13932
rect 8803 13892 9496 13920
rect 8803 13889 8815 13892
rect 8757 13883 8815 13889
rect 9490 13880 9496 13892
rect 9548 13920 9554 13932
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 9548 13892 10425 13920
rect 9548 13880 9554 13892
rect 10413 13889 10425 13892
rect 10459 13920 10471 13923
rect 11238 13920 11244 13932
rect 10459 13892 11244 13920
rect 10459 13889 10471 13892
rect 10413 13883 10471 13889
rect 11238 13880 11244 13892
rect 11296 13920 11302 13932
rect 11296 13892 12204 13920
rect 11296 13880 11302 13892
rect 5399 13824 6040 13852
rect 6089 13855 6147 13861
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 6089 13821 6101 13855
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 5258 13784 5264 13796
rect 4724 13756 5264 13784
rect 5258 13744 5264 13756
rect 5316 13744 5322 13796
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6104 13784 6132 13815
rect 6914 13812 6920 13864
rect 6972 13812 6978 13864
rect 7006 13812 7012 13864
rect 7064 13812 7070 13864
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8662 13852 8668 13864
rect 7883 13824 8668 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 8662 13812 8668 13824
rect 8720 13812 8726 13864
rect 8846 13812 8852 13864
rect 8904 13852 8910 13864
rect 10226 13852 10232 13864
rect 8904 13824 10232 13852
rect 8904 13812 8910 13824
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10594 13852 10600 13864
rect 10367 13824 10600 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10778 13812 10784 13864
rect 10836 13812 10842 13864
rect 11790 13852 11796 13864
rect 11026 13824 11796 13852
rect 11026 13784 11054 13824
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 12176 13861 12204 13892
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13821 12127 13855
rect 12069 13815 12127 13821
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13852 12219 13855
rect 12805 13855 12863 13861
rect 12805 13852 12817 13855
rect 12207 13824 12817 13852
rect 12207 13821 12219 13824
rect 12161 13815 12219 13821
rect 12805 13821 12817 13824
rect 12851 13821 12863 13855
rect 12805 13815 12863 13821
rect 5592 13756 11054 13784
rect 12084 13784 12112 13815
rect 12894 13812 12900 13864
rect 12952 13852 12958 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12952 13824 13001 13852
rect 12952 13812 12958 13824
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 12989 13815 13047 13821
rect 13262 13812 13268 13864
rect 13320 13812 13326 13864
rect 13541 13855 13599 13861
rect 13541 13821 13553 13855
rect 13587 13821 13599 13855
rect 13541 13815 13599 13821
rect 12710 13784 12716 13796
rect 12084 13756 12716 13784
rect 5592 13744 5598 13756
rect 12710 13744 12716 13756
rect 12768 13784 12774 13796
rect 13556 13784 13584 13815
rect 14090 13812 14096 13864
rect 14148 13812 14154 13864
rect 12768 13756 13584 13784
rect 12768 13744 12774 13756
rect 6454 13676 6460 13728
rect 6512 13676 6518 13728
rect 7377 13719 7435 13725
rect 7377 13685 7389 13719
rect 7423 13716 7435 13719
rect 7466 13716 7472 13728
rect 7423 13688 7472 13716
rect 7423 13685 7435 13688
rect 7377 13679 7435 13685
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 8205 13719 8263 13725
rect 8205 13685 8217 13719
rect 8251 13716 8263 13719
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 8251 13688 8401 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8389 13685 8401 13688
rect 8435 13685 8447 13719
rect 8389 13679 8447 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 10594 13716 10600 13728
rect 8720 13688 10600 13716
rect 8720 13676 8726 13688
rect 10594 13676 10600 13688
rect 10652 13716 10658 13728
rect 11238 13716 11244 13728
rect 10652 13688 11244 13716
rect 10652 13676 10658 13688
rect 11238 13676 11244 13688
rect 11296 13716 11302 13728
rect 11609 13719 11667 13725
rect 11609 13716 11621 13719
rect 11296 13688 11621 13716
rect 11296 13676 11302 13688
rect 11609 13685 11621 13688
rect 11655 13685 11667 13719
rect 11609 13679 11667 13685
rect 12529 13719 12587 13725
rect 12529 13685 12541 13719
rect 12575 13716 12587 13719
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12575 13688 12633 13716
rect 12575 13685 12587 13688
rect 12529 13679 12587 13685
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 12621 13679 12679 13685
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 13081 13719 13139 13725
rect 13081 13716 13093 13719
rect 13044 13688 13093 13716
rect 13044 13676 13050 13688
rect 13081 13685 13093 13688
rect 13127 13685 13139 13719
rect 13081 13679 13139 13685
rect 13633 13719 13691 13725
rect 13633 13685 13645 13719
rect 13679 13716 13691 13719
rect 13814 13716 13820 13728
rect 13679 13688 13820 13716
rect 13679 13685 13691 13688
rect 13633 13679 13691 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 5123 13484 5181 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 7377 13515 7435 13521
rect 7377 13481 7389 13515
rect 7423 13512 7435 13515
rect 7466 13512 7472 13524
rect 7423 13484 7472 13512
rect 7423 13481 7435 13484
rect 7377 13475 7435 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 10962 13512 10968 13524
rect 7576 13484 10968 13512
rect 3234 13404 3240 13456
rect 3292 13444 3298 13456
rect 3292 13416 4108 13444
rect 3292 13404 3298 13416
rect 4080 13385 4108 13416
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 6058 13447 6116 13453
rect 6058 13444 6070 13447
rect 5776 13416 6070 13444
rect 5776 13404 5782 13416
rect 6058 13413 6070 13416
rect 6104 13413 6116 13447
rect 6058 13407 6116 13413
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7576 13444 7604 13484
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11238 13472 11244 13524
rect 11296 13512 11302 13524
rect 12894 13512 12900 13524
rect 11296 13484 12900 13512
rect 11296 13472 11302 13484
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 6972 13416 7604 13444
rect 6972 13404 6978 13416
rect 8846 13404 8852 13456
rect 8904 13444 8910 13456
rect 10042 13444 10048 13456
rect 8904 13416 10048 13444
rect 8904 13404 8910 13416
rect 10042 13404 10048 13416
rect 10100 13444 10106 13456
rect 10689 13447 10747 13453
rect 10689 13444 10701 13447
rect 10100 13416 10701 13444
rect 10100 13404 10106 13416
rect 10689 13413 10701 13416
rect 10735 13413 10747 13447
rect 10689 13407 10747 13413
rect 15013 13447 15071 13453
rect 15013 13413 15025 13447
rect 15059 13444 15071 13447
rect 15102 13444 15108 13456
rect 15059 13416 15108 13444
rect 15059 13413 15071 13416
rect 15013 13407 15071 13413
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 3809 13379 3867 13385
rect 3809 13345 3821 13379
rect 3855 13376 3867 13379
rect 4065 13379 4123 13385
rect 3855 13348 4016 13376
rect 3855 13345 3867 13348
rect 3809 13339 3867 13345
rect 3988 13308 4016 13348
rect 4065 13345 4077 13379
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 5166 13376 5172 13388
rect 4755 13348 5172 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5353 13379 5411 13385
rect 5353 13376 5365 13379
rect 5316 13348 5365 13376
rect 5316 13336 5322 13348
rect 5353 13345 5365 13348
rect 5399 13345 5411 13379
rect 5353 13339 5411 13345
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 5810 13336 5816 13388
rect 5868 13336 5874 13388
rect 7650 13336 7656 13388
rect 7708 13336 7714 13388
rect 7745 13379 7803 13385
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 8662 13376 8668 13388
rect 7791 13348 8668 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9398 13385 9404 13388
rect 9392 13339 9404 13385
rect 9398 13336 9404 13339
rect 9456 13336 9462 13388
rect 10597 13379 10655 13385
rect 10597 13376 10609 13379
rect 10520 13348 10609 13376
rect 4433 13311 4491 13317
rect 4433 13308 4445 13311
rect 3988 13280 4445 13308
rect 4433 13277 4445 13280
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 7668 13308 7696 13336
rect 8757 13311 8815 13317
rect 8757 13308 8769 13311
rect 7668 13280 8769 13308
rect 4617 13271 4675 13277
rect 8757 13277 8769 13280
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 4632 13240 4660 13271
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 4982 13240 4988 13252
rect 4632 13212 4988 13240
rect 4982 13200 4988 13212
rect 5040 13240 5046 13252
rect 8938 13240 8944 13252
rect 5040 13212 5488 13240
rect 5040 13200 5046 13212
rect 2685 13175 2743 13181
rect 2685 13141 2697 13175
rect 2731 13172 2743 13175
rect 4798 13172 4804 13184
rect 2731 13144 4804 13172
rect 2731 13141 2743 13144
rect 2685 13135 2743 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 4890 13132 4896 13184
rect 4948 13172 4954 13184
rect 5353 13175 5411 13181
rect 5353 13172 5365 13175
rect 4948 13144 5365 13172
rect 4948 13132 4954 13144
rect 5353 13141 5365 13144
rect 5399 13141 5411 13175
rect 5460 13172 5488 13212
rect 6840 13212 8944 13240
rect 6840 13172 6868 13212
rect 8938 13200 8944 13212
rect 8996 13200 9002 13252
rect 10520 13249 10548 13348
rect 10597 13345 10609 13348
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13376 11575 13379
rect 11882 13376 11888 13388
rect 11563 13348 11888 13376
rect 11563 13345 11575 13348
rect 11517 13339 11575 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12986 13336 12992 13388
rect 13044 13336 13050 13388
rect 13170 13336 13176 13388
rect 13228 13376 13234 13388
rect 13633 13379 13691 13385
rect 13633 13376 13645 13379
rect 13228 13348 13645 13376
rect 13228 13336 13234 13348
rect 13633 13345 13645 13348
rect 13679 13345 13691 13379
rect 13633 13339 13691 13345
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 13136 13280 13277 13308
rect 13136 13268 13142 13280
rect 13265 13277 13277 13280
rect 13311 13308 13323 13311
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 13311 13280 13369 13308
rect 13311 13277 13323 13280
rect 13265 13271 13323 13277
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 10505 13243 10563 13249
rect 10505 13209 10517 13243
rect 10551 13209 10563 13243
rect 10505 13203 10563 13209
rect 5460 13144 6868 13172
rect 5353 13135 5411 13141
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 6972 13144 7205 13172
rect 6972 13132 6978 13144
rect 7193 13141 7205 13144
rect 7239 13141 7251 13175
rect 7193 13135 7251 13141
rect 7558 13132 7564 13184
rect 7616 13132 7622 13184
rect 8846 13132 8852 13184
rect 8904 13132 8910 13184
rect 9030 13132 9036 13184
rect 9088 13132 9094 13184
rect 11422 13132 11428 13184
rect 11480 13132 11486 13184
rect 11514 13132 11520 13184
rect 11572 13172 11578 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11572 13144 11897 13172
rect 11572 13132 11578 13144
rect 11885 13141 11897 13144
rect 11931 13172 11943 13175
rect 13078 13172 13084 13184
rect 11931 13144 13084 13172
rect 11931 13141 11943 13144
rect 11885 13135 11943 13141
rect 13078 13132 13084 13144
rect 13136 13132 13142 13184
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 4890 12928 4896 12980
rect 4948 12928 4954 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5776 12940 5825 12968
rect 5776 12928 5782 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 6270 12928 6276 12980
rect 6328 12968 6334 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 6328 12940 6837 12968
rect 6328 12928 6334 12940
rect 6825 12937 6837 12940
rect 6871 12968 6883 12971
rect 7190 12968 7196 12980
rect 6871 12940 7196 12968
rect 6871 12937 6883 12940
rect 6825 12931 6883 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 9398 12928 9404 12980
rect 9456 12968 9462 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9456 12940 9873 12968
rect 9456 12928 9462 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 13262 12968 13268 12980
rect 11931 12940 13268 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 4614 12832 4620 12844
rect 4356 12804 4620 12832
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 4356 12773 4384 12804
rect 4614 12792 4620 12804
rect 4672 12832 4678 12844
rect 4908 12832 4936 12928
rect 7466 12860 7472 12912
rect 7524 12900 7530 12912
rect 8665 12903 8723 12909
rect 8665 12900 8677 12903
rect 7524 12872 8677 12900
rect 7524 12860 7530 12872
rect 8665 12869 8677 12872
rect 8711 12869 8723 12903
rect 8665 12863 8723 12869
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 8996 12872 12112 12900
rect 8996 12860 9002 12872
rect 6089 12835 6147 12841
rect 6089 12832 6101 12835
rect 4672 12804 4936 12832
rect 5506 12804 6101 12832
rect 4672 12792 4678 12804
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 4706 12764 4712 12776
rect 4580 12736 4712 12764
rect 4580 12724 4586 12736
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 4798 12724 4804 12776
rect 4856 12724 4862 12776
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5506 12764 5534 12804
rect 6089 12801 6101 12804
rect 6135 12801 6147 12835
rect 6089 12795 6147 12801
rect 6454 12792 6460 12844
rect 6512 12792 6518 12844
rect 8570 12832 8576 12844
rect 6840 12804 8576 12832
rect 5224 12736 5534 12764
rect 5997 12767 6055 12773
rect 5224 12724 5230 12736
rect 5997 12733 6009 12767
rect 6043 12764 6055 12767
rect 6362 12764 6368 12776
rect 6043 12736 6368 12764
rect 6043 12733 6055 12736
rect 5997 12727 6055 12733
rect 6362 12724 6368 12736
rect 6420 12764 6426 12776
rect 6840 12764 6868 12804
rect 8570 12792 8576 12804
rect 8628 12792 8634 12844
rect 9030 12792 9036 12844
rect 9088 12832 9094 12844
rect 9217 12835 9275 12841
rect 9217 12832 9229 12835
rect 9088 12804 9229 12832
rect 9088 12792 9094 12804
rect 9217 12801 9229 12804
rect 9263 12801 9275 12835
rect 9217 12795 9275 12801
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9548 12804 9597 12832
rect 9548 12792 9554 12804
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 11422 12832 11428 12844
rect 10836 12804 11428 12832
rect 10836 12792 10842 12804
rect 11422 12792 11428 12804
rect 11480 12832 11486 12844
rect 12084 12841 12112 12872
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11480 12804 11529 12832
rect 11480 12792 11486 12804
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12832 12495 12835
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12483 12804 12817 12832
rect 12483 12801 12495 12804
rect 12437 12795 12495 12801
rect 12805 12801 12817 12804
rect 12851 12832 12863 12835
rect 13817 12835 13875 12841
rect 13817 12832 13829 12835
rect 12851 12804 13829 12832
rect 12851 12801 12863 12804
rect 12805 12795 12863 12801
rect 13817 12801 13829 12804
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 6420 12736 6868 12764
rect 6420 12724 6426 12736
rect 6914 12724 6920 12776
rect 6972 12724 6978 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10410 12764 10416 12776
rect 9723 12736 10416 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 11701 12767 11759 12773
rect 11701 12733 11713 12767
rect 11747 12764 11759 12767
rect 11882 12764 11888 12776
rect 11747 12736 11888 12764
rect 11747 12733 11759 12736
rect 11701 12727 11759 12733
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 12342 12724 12348 12776
rect 12400 12724 12406 12776
rect 12710 12724 12716 12776
rect 12768 12764 12774 12776
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12768 12736 13001 12764
rect 12768 12724 12774 12736
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13078 12724 13084 12776
rect 13136 12764 13142 12776
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 13136 12736 13185 12764
rect 13136 12724 13142 12736
rect 13173 12733 13185 12736
rect 13219 12764 13231 12767
rect 13262 12764 13268 12776
rect 13219 12736 13268 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13906 12724 13912 12776
rect 13964 12764 13970 12776
rect 15102 12764 15108 12776
rect 13964 12736 15108 12764
rect 13964 12724 13970 12736
rect 15102 12724 15108 12736
rect 15160 12724 15166 12776
rect 4430 12656 4436 12708
rect 4488 12696 4494 12708
rect 5350 12696 5356 12708
rect 4488 12668 5356 12696
rect 4488 12656 4494 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 8352 12668 8401 12696
rect 8352 12656 8358 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 8389 12659 8447 12665
rect 11977 12699 12035 12705
rect 11977 12665 11989 12699
rect 12023 12696 12035 12699
rect 12158 12696 12164 12708
rect 12023 12668 12164 12696
rect 12023 12665 12035 12668
rect 11977 12659 12035 12665
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 4706 12588 4712 12640
rect 4764 12588 4770 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7558 12628 7564 12640
rect 7064 12600 7564 12628
rect 7064 12588 7070 12600
rect 7558 12588 7564 12600
rect 7616 12588 7622 12640
rect 8849 12631 8907 12637
rect 8849 12597 8861 12631
rect 8895 12628 8907 12631
rect 9030 12628 9036 12640
rect 8895 12600 9036 12628
rect 8895 12597 8907 12600
rect 8849 12591 8907 12597
rect 9030 12588 9036 12600
rect 9088 12588 9094 12640
rect 12618 12588 12624 12640
rect 12676 12588 12682 12640
rect 13541 12631 13599 12637
rect 13541 12597 13553 12631
rect 13587 12628 13599 12631
rect 13722 12628 13728 12640
rect 13587 12600 13728 12628
rect 13587 12597 13599 12600
rect 13541 12591 13599 12597
rect 13722 12588 13728 12600
rect 13780 12588 13786 12640
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 8110 12424 8116 12436
rect 4663 12396 8116 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8662 12424 8668 12436
rect 8444 12396 8668 12424
rect 8444 12384 8450 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11422 12424 11428 12436
rect 11379 12396 11428 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11422 12384 11428 12396
rect 11480 12384 11486 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 11882 12424 11888 12436
rect 11747 12396 11888 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 4249 12359 4307 12365
rect 4249 12325 4261 12359
rect 4295 12356 4307 12359
rect 4709 12359 4767 12365
rect 4709 12356 4721 12359
rect 4295 12328 4721 12356
rect 4295 12325 4307 12328
rect 4249 12319 4307 12325
rect 4709 12325 4721 12328
rect 4755 12325 4767 12359
rect 4709 12319 4767 12325
rect 7101 12359 7159 12365
rect 7101 12325 7113 12359
rect 7147 12356 7159 12359
rect 7147 12328 7328 12356
rect 7147 12325 7159 12328
rect 7101 12319 7159 12325
rect 7300 12300 7328 12328
rect 7466 12316 7472 12368
rect 7524 12316 7530 12368
rect 8404 12356 8432 12384
rect 8036 12328 8432 12356
rect 11241 12359 11299 12365
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 4154 12297 4160 12300
rect 3973 12291 4031 12297
rect 3973 12288 3985 12291
rect 3660 12260 3985 12288
rect 3660 12248 3666 12260
rect 3973 12257 3985 12260
rect 4019 12257 4031 12291
rect 3973 12251 4031 12257
rect 4121 12291 4160 12297
rect 4121 12257 4133 12291
rect 4121 12251 4160 12257
rect 4154 12248 4160 12251
rect 4212 12248 4218 12300
rect 4338 12248 4344 12300
rect 4396 12248 4402 12300
rect 4438 12291 4496 12297
rect 4438 12257 4450 12291
rect 4484 12288 4496 12291
rect 4484 12260 4568 12288
rect 4484 12257 4496 12260
rect 4438 12251 4496 12257
rect 4540 12232 4568 12260
rect 4798 12248 4804 12300
rect 4856 12288 4862 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4856 12260 4905 12288
rect 4856 12248 4862 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 4893 12251 4951 12257
rect 5169 12291 5227 12297
rect 5169 12257 5181 12291
rect 5215 12257 5227 12291
rect 5169 12251 5227 12257
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 5184 12220 5212 12251
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5626 12288 5632 12300
rect 5408 12260 5632 12288
rect 5408 12248 5414 12260
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 6871 12260 6960 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 4580 12192 5212 12220
rect 4580 12180 4586 12192
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 5442 12084 5448 12096
rect 3835 12056 5448 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6546 12044 6552 12096
rect 6604 12084 6610 12096
rect 6932 12084 6960 12260
rect 7006 12248 7012 12300
rect 7064 12248 7070 12300
rect 7190 12248 7196 12300
rect 7248 12248 7254 12300
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7742 12288 7748 12300
rect 7699 12260 7748 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 8036 12297 8064 12328
rect 11241 12325 11253 12359
rect 11287 12356 11299 12359
rect 12618 12356 12624 12368
rect 11287 12328 12624 12356
rect 11287 12325 11299 12328
rect 11241 12319 11299 12325
rect 12618 12316 12624 12328
rect 12676 12316 12682 12368
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12257 8079 12291
rect 8021 12251 8079 12257
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7616 12192 7849 12220
rect 7616 12180 7622 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 7926 12180 7932 12232
rect 7984 12180 7990 12232
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8312 12220 8340 12251
rect 8386 12248 8392 12300
rect 8444 12248 8450 12300
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 8536 12260 8585 12288
rect 8536 12248 8542 12260
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12257 8723 12291
rect 8665 12251 8723 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12257 8815 12291
rect 8757 12251 8815 12257
rect 8168 12192 8340 12220
rect 8168 12180 8174 12192
rect 7377 12155 7435 12161
rect 7377 12121 7389 12155
rect 7423 12152 7435 12155
rect 8294 12152 8300 12164
rect 7423 12124 8300 12152
rect 7423 12121 7435 12124
rect 7377 12115 7435 12121
rect 8294 12112 8300 12124
rect 8352 12152 8358 12164
rect 8680 12152 8708 12251
rect 8352 12124 8708 12152
rect 8352 12112 8358 12124
rect 7742 12084 7748 12096
rect 6604 12056 7748 12084
rect 6604 12044 6610 12056
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8772 12084 8800 12251
rect 11790 12248 11796 12300
rect 11848 12248 11854 12300
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 8941 12155 8999 12161
rect 8941 12121 8953 12155
rect 8987 12152 8999 12155
rect 11054 12152 11060 12164
rect 8987 12124 11060 12152
rect 8987 12121 8999 12124
rect 8941 12115 8999 12121
rect 11054 12112 11060 12124
rect 11112 12152 11118 12164
rect 11164 12152 11192 12183
rect 11112 12124 11192 12152
rect 11112 12112 11118 12124
rect 8260 12056 8800 12084
rect 8260 12044 8266 12056
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 13044 12056 13093 12084
rect 13044 12044 13050 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 4522 11880 4528 11892
rect 4387 11852 4528 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 5074 11840 5080 11892
rect 5132 11880 5138 11892
rect 5132 11852 5304 11880
rect 5132 11840 5138 11852
rect 4801 11815 4859 11821
rect 4801 11781 4813 11815
rect 4847 11812 4859 11815
rect 5169 11815 5227 11821
rect 5169 11812 5181 11815
rect 4847 11784 5181 11812
rect 4847 11781 4859 11784
rect 4801 11775 4859 11781
rect 5169 11781 5181 11784
rect 5215 11781 5227 11815
rect 5276 11812 5304 11852
rect 7374 11840 7380 11892
rect 7432 11840 7438 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8481 11883 8539 11889
rect 8481 11880 8493 11883
rect 8444 11852 8493 11880
rect 8444 11840 8450 11852
rect 8481 11849 8493 11852
rect 8527 11849 8539 11883
rect 8481 11843 8539 11849
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8628 11852 11744 11880
rect 8628 11840 8634 11852
rect 11146 11812 11152 11824
rect 5276 11784 10916 11812
rect 5169 11775 5227 11781
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 4212 11716 4568 11744
rect 4212 11704 4218 11716
rect 4540 11688 4568 11716
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 10888 11753 10916 11784
rect 10980 11784 11152 11812
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4764 11716 4905 11744
rect 4764 11704 4770 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 10321 11747 10379 11753
rect 10321 11744 10333 11747
rect 4893 11707 4951 11713
rect 8864 11716 10333 11744
rect 4249 11679 4307 11685
rect 4249 11645 4261 11679
rect 4295 11676 4307 11679
rect 4430 11676 4436 11688
rect 4295 11648 4436 11676
rect 4295 11645 4307 11648
rect 4249 11639 4307 11645
rect 4430 11636 4436 11648
rect 4488 11636 4494 11688
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 8754 11636 8760 11688
rect 8812 11636 8818 11688
rect 8864 11685 8892 11716
rect 10321 11713 10333 11716
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11645 8999 11679
rect 8941 11639 8999 11645
rect 6089 11611 6147 11617
rect 6089 11577 6101 11611
rect 6135 11608 6147 11611
rect 7650 11608 7656 11620
rect 6135 11580 7656 11608
rect 6135 11577 6147 11580
rect 6089 11571 6147 11577
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 8478 11608 8484 11620
rect 7852 11580 8484 11608
rect 5353 11543 5411 11549
rect 5353 11509 5365 11543
rect 5399 11540 5411 11543
rect 7852 11540 7880 11580
rect 8478 11568 8484 11580
rect 8536 11608 8542 11620
rect 8956 11608 8984 11639
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9125 11679 9183 11685
rect 9125 11676 9137 11679
rect 9088 11648 9137 11676
rect 9088 11636 9094 11648
rect 9125 11645 9137 11648
rect 9171 11645 9183 11679
rect 9125 11639 9183 11645
rect 9582 11636 9588 11688
rect 9640 11636 9646 11688
rect 9766 11676 9772 11688
rect 9692 11648 9772 11676
rect 8536 11580 8984 11608
rect 9692 11608 9720 11648
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 9858 11636 9864 11688
rect 9916 11636 9922 11688
rect 9953 11679 10011 11685
rect 9953 11645 9965 11679
rect 9999 11676 10011 11679
rect 10042 11676 10048 11688
rect 9999 11648 10048 11676
rect 9999 11645 10011 11648
rect 9953 11639 10011 11645
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 10134 11636 10140 11688
rect 10192 11636 10198 11688
rect 10686 11636 10692 11688
rect 10744 11676 10750 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10744 11648 10793 11676
rect 10744 11636 10750 11648
rect 10781 11645 10793 11648
rect 10827 11676 10839 11679
rect 10980 11676 11008 11784
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 11057 11747 11115 11753
rect 11057 11713 11069 11747
rect 11103 11744 11115 11747
rect 11422 11744 11428 11756
rect 11103 11716 11428 11744
rect 11103 11713 11115 11716
rect 11057 11707 11115 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 11716 11685 11744 11852
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12621 11883 12679 11889
rect 12621 11880 12633 11883
rect 12400 11852 12633 11880
rect 12400 11840 12406 11852
rect 12621 11849 12633 11852
rect 12667 11849 12679 11883
rect 12621 11843 12679 11849
rect 12710 11840 12716 11892
rect 12768 11840 12774 11892
rect 11808 11784 13584 11812
rect 11333 11679 11391 11685
rect 11333 11676 11345 11679
rect 10827 11648 11008 11676
rect 11072 11648 11345 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 11072 11620 11100 11648
rect 11333 11645 11345 11648
rect 11379 11645 11391 11679
rect 11333 11639 11391 11645
rect 11701 11679 11759 11685
rect 11701 11645 11713 11679
rect 11747 11645 11759 11679
rect 11701 11639 11759 11645
rect 10502 11608 10508 11620
rect 9692 11580 10508 11608
rect 8536 11568 8542 11580
rect 10502 11568 10508 11580
rect 10560 11568 10566 11620
rect 11054 11568 11060 11620
rect 11112 11568 11118 11620
rect 11146 11568 11152 11620
rect 11204 11608 11210 11620
rect 11808 11608 11836 11784
rect 12529 11747 12587 11753
rect 12529 11744 12541 11747
rect 12268 11716 12541 11744
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 11204 11580 11836 11608
rect 11204 11568 11210 11580
rect 5399 11512 7880 11540
rect 5399 11509 5411 11512
rect 5353 11503 5411 11509
rect 7926 11500 7932 11552
rect 7984 11540 7990 11552
rect 8570 11540 8576 11552
rect 7984 11512 8576 11540
rect 7984 11500 7990 11512
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10594 11540 10600 11552
rect 10459 11512 10600 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 10928 11512 11529 11540
rect 10928 11500 10934 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 11882 11540 11888 11552
rect 11839 11512 11888 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12268 11549 12296 11716
rect 12529 11713 12541 11716
rect 12575 11713 12587 11747
rect 12529 11707 12587 11713
rect 12805 11679 12863 11685
rect 12805 11645 12817 11679
rect 12851 11676 12863 11679
rect 13262 11676 13268 11688
rect 12851 11648 13268 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 13262 11636 13268 11648
rect 13320 11636 13326 11688
rect 13556 11685 13584 11784
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11645 13599 11679
rect 13541 11639 13599 11645
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 12124 11512 12265 11540
rect 12124 11500 12130 11512
rect 12253 11509 12265 11512
rect 12299 11509 12311 11543
rect 12253 11503 12311 11509
rect 12802 11500 12808 11552
rect 12860 11540 12866 11552
rect 13633 11543 13691 11549
rect 13633 11540 13645 11543
rect 12860 11512 13645 11540
rect 12860 11500 12866 11512
rect 13633 11509 13645 11512
rect 13679 11509 13691 11543
rect 13633 11503 13691 11509
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8202 11336 8208 11348
rect 7791 11308 8208 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8202 11296 8208 11308
rect 8260 11296 8266 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 8754 11336 8760 11348
rect 8527 11308 8760 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 8754 11296 8760 11308
rect 8812 11296 8818 11348
rect 9582 11296 9588 11348
rect 9640 11296 9646 11348
rect 10042 11296 10048 11348
rect 10100 11296 10106 11348
rect 11054 11336 11060 11348
rect 10428 11308 11060 11336
rect 6080 11271 6138 11277
rect 6080 11237 6092 11271
rect 6126 11268 6138 11271
rect 6270 11268 6276 11280
rect 6126 11240 6276 11268
rect 6126 11237 6138 11240
rect 6080 11231 6138 11237
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 8849 11271 8907 11277
rect 8628 11240 8800 11268
rect 8628 11228 8634 11240
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 5718 11200 5724 11212
rect 5399 11172 5724 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 5184 11132 5212 11163
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 5810 11160 5816 11212
rect 5868 11160 5874 11212
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 7285 11203 7343 11209
rect 7285 11200 7297 11203
rect 6972 11172 7297 11200
rect 6972 11160 6978 11172
rect 7285 11169 7297 11172
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11169 7895 11203
rect 7837 11163 7895 11169
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 5534 11132 5540 11144
rect 5184 11104 5540 11132
rect 5534 11092 5540 11104
rect 5592 11092 5598 11144
rect 7852 11132 7880 11163
rect 7208 11104 7880 11132
rect 5350 10956 5356 11008
rect 5408 10956 5414 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 7208 11005 7236 11104
rect 8036 11064 8064 11163
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8772 11209 8800 11240
rect 8849 11237 8861 11271
rect 8895 11268 8907 11271
rect 10060 11268 10088 11296
rect 10428 11277 10456 11308
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 11701 11339 11759 11345
rect 11701 11305 11713 11339
rect 11747 11336 11759 11339
rect 11882 11336 11888 11348
rect 11747 11308 11888 11336
rect 11747 11305 11759 11308
rect 11701 11299 11759 11305
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13228 11308 13277 11336
rect 13228 11296 13234 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 8895 11240 10088 11268
rect 10413 11271 10471 11277
rect 8895 11237 8907 11240
rect 8849 11231 8907 11237
rect 10413 11237 10425 11271
rect 10459 11237 10471 11271
rect 10413 11231 10471 11237
rect 11422 11228 11428 11280
rect 11480 11268 11486 11280
rect 11480 11240 12756 11268
rect 11480 11228 11486 11240
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8996 11172 9045 11200
rect 8996 11160 9002 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 9766 11160 9772 11212
rect 9824 11160 9830 11212
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 10045 11203 10103 11209
rect 10045 11169 10057 11203
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 10226 11200 10232 11212
rect 10183 11172 10232 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 9876 11132 9904 11160
rect 9364 11104 9904 11132
rect 10060 11132 10088 11163
rect 10226 11160 10232 11172
rect 10284 11160 10290 11212
rect 10962 11160 10968 11212
rect 11020 11160 11026 11212
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 11793 11203 11851 11209
rect 11793 11169 11805 11203
rect 11839 11169 11851 11203
rect 11793 11163 11851 11169
rect 12529 11203 12587 11209
rect 12529 11169 12541 11203
rect 12575 11200 12587 11203
rect 12618 11200 12624 11212
rect 12575 11172 12624 11200
rect 12575 11169 12587 11172
rect 12529 11163 12587 11169
rect 10060 11104 11054 11132
rect 9364 11092 9370 11104
rect 10686 11064 10692 11076
rect 8036 11036 10692 11064
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 11026 11064 11054 11104
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 11808 11132 11836 11163
rect 12618 11160 12624 11172
rect 12676 11160 12682 11212
rect 12728 11209 12756 11240
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11169 12771 11203
rect 12713 11163 12771 11169
rect 12802 11160 12808 11212
rect 12860 11160 12866 11212
rect 13081 11203 13139 11209
rect 13081 11169 13093 11203
rect 13127 11200 13139 11203
rect 13906 11200 13912 11212
rect 13127 11172 13912 11200
rect 13127 11169 13139 11172
rect 13081 11163 13139 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 12434 11132 12440 11144
rect 11808 11104 12440 11132
rect 12434 11092 12440 11104
rect 12492 11092 12498 11144
rect 12894 11092 12900 11144
rect 12952 11092 12958 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 13044 11104 13369 11132
rect 13044 11092 13050 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13630 11092 13636 11144
rect 13688 11092 13694 11144
rect 11882 11064 11888 11076
rect 11026 11036 11888 11064
rect 11882 11024 11888 11036
rect 11940 11024 11946 11076
rect 11974 11024 11980 11076
rect 12032 11064 12038 11076
rect 12032 11036 12388 11064
rect 12032 11024 12038 11036
rect 7193 10999 7251 11005
rect 7193 10996 7205 10999
rect 5684 10968 7205 10996
rect 5684 10956 5690 10968
rect 7193 10965 7205 10968
rect 7239 10965 7251 10999
rect 7193 10959 7251 10965
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 7377 10999 7435 11005
rect 7377 10996 7389 10999
rect 7340 10968 7389 10996
rect 7340 10956 7346 10968
rect 7377 10965 7389 10968
rect 7423 10965 7435 10999
rect 7377 10959 7435 10965
rect 7926 10956 7932 11008
rect 7984 10956 7990 11008
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10996 10379 10999
rect 10594 10996 10600 11008
rect 10367 10968 10600 10996
rect 10367 10965 10379 10968
rect 10321 10959 10379 10965
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 11057 10999 11115 11005
rect 11057 10965 11069 10999
rect 11103 10996 11115 10999
rect 11238 10996 11244 11008
rect 11103 10968 11244 10996
rect 11103 10965 11115 10968
rect 11057 10959 11115 10965
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 12158 10956 12164 11008
rect 12216 10956 12222 11008
rect 12360 10996 12388 11036
rect 12544 11036 13400 11064
rect 12544 10996 12572 11036
rect 12360 10968 12572 10996
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13170 10996 13176 11008
rect 12952 10968 13176 10996
rect 12952 10956 12958 10968
rect 13170 10956 13176 10968
rect 13228 10956 13234 11008
rect 13372 10996 13400 11036
rect 13630 10996 13636 11008
rect 13372 10968 13636 10996
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 14921 10999 14979 11005
rect 14921 10965 14933 10999
rect 14967 10996 14979 10999
rect 15102 10996 15108 11008
rect 14967 10968 15108 10996
rect 14967 10965 14979 10968
rect 14921 10959 14979 10965
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 6181 10795 6239 10801
rect 4632 10764 5488 10792
rect 4632 10665 4660 10764
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 5460 10724 5488 10764
rect 6181 10761 6193 10795
rect 6227 10792 6239 10795
rect 6270 10792 6276 10804
rect 6227 10764 6276 10792
rect 6227 10761 6239 10764
rect 6181 10755 6239 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 7374 10792 7380 10804
rect 6503 10764 7380 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 7374 10752 7380 10764
rect 7432 10792 7438 10804
rect 9582 10792 9588 10804
rect 7432 10764 9588 10792
rect 7432 10752 7438 10764
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 12250 10792 12256 10804
rect 11664 10764 12256 10792
rect 11664 10752 11670 10764
rect 12250 10752 12256 10764
rect 12308 10792 12314 10804
rect 12526 10792 12532 10804
rect 12308 10764 12532 10792
rect 12308 10752 12314 10764
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12768 10764 12817 10792
rect 12768 10752 12774 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 12989 10795 13047 10801
rect 12989 10792 13001 10795
rect 12952 10764 13001 10792
rect 12952 10752 12958 10764
rect 12989 10761 13001 10764
rect 13035 10792 13047 10795
rect 13035 10764 14412 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 5810 10724 5816 10736
rect 5316 10696 5396 10724
rect 5460 10696 5816 10724
rect 5316 10684 5322 10696
rect 5368 10665 5396 10696
rect 5810 10684 5816 10696
rect 5868 10684 5874 10736
rect 6549 10727 6607 10733
rect 6549 10693 6561 10727
rect 6595 10693 6607 10727
rect 6549 10687 6607 10693
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6564 10656 6592 10687
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9677 10727 9735 10733
rect 9677 10724 9689 10727
rect 9272 10696 9689 10724
rect 9272 10684 9278 10696
rect 9677 10693 9689 10696
rect 9723 10693 9735 10727
rect 14277 10727 14335 10733
rect 14277 10724 14289 10727
rect 9677 10687 9735 10693
rect 11900 10696 14289 10724
rect 5767 10628 6592 10656
rect 6641 10659 6699 10665
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 7926 10656 7932 10668
rect 6687 10628 7932 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 8444 10628 9321 10656
rect 8444 10616 8450 10628
rect 9309 10625 9321 10628
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 10962 10616 10968 10668
rect 11020 10656 11026 10668
rect 11609 10659 11667 10665
rect 11609 10656 11621 10659
rect 11020 10628 11621 10656
rect 11020 10616 11026 10628
rect 11609 10625 11621 10628
rect 11655 10625 11667 10659
rect 11609 10619 11667 10625
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 5224 10560 5457 10588
rect 5224 10548 5230 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 5445 10551 5503 10557
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5813 10591 5871 10597
rect 5813 10557 5825 10591
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6365 10591 6423 10597
rect 6365 10588 6377 10591
rect 6043 10560 6377 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6365 10557 6377 10560
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 4372 10523 4430 10529
rect 4372 10489 4384 10523
rect 4418 10520 4430 10523
rect 4614 10520 4620 10532
rect 4418 10492 4620 10520
rect 4418 10489 4430 10492
rect 4372 10483 4430 10489
rect 4614 10480 4620 10492
rect 4672 10480 4678 10532
rect 5350 10480 5356 10532
rect 5408 10520 5414 10532
rect 5644 10520 5672 10551
rect 5408 10492 5672 10520
rect 5408 10480 5414 10492
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 5828 10520 5856 10551
rect 5776 10492 5856 10520
rect 5776 10480 5782 10492
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 4522 10452 4528 10464
rect 3283 10424 4528 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4890 10452 4896 10464
rect 4755 10424 4896 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6012 10452 6040 10551
rect 8938 10548 8944 10600
rect 8996 10588 9002 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8996 10560 9137 10588
rect 8996 10548 9002 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9140 10520 9168 10551
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 10134 10588 10140 10600
rect 9508 10560 10140 10588
rect 9508 10529 9536 10560
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11204 10560 11529 10588
rect 11204 10548 11210 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11900 10588 11928 10696
rect 14277 10693 14289 10696
rect 14323 10693 14335 10727
rect 14277 10687 14335 10693
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10656 12035 10659
rect 12158 10656 12164 10668
rect 12023 10628 12164 10656
rect 12023 10625 12035 10628
rect 11977 10619 12035 10625
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11900 10560 12081 10588
rect 11517 10551 11575 10557
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12250 10548 12256 10600
rect 12308 10548 12314 10600
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 9493 10523 9551 10529
rect 9493 10520 9505 10523
rect 9140 10492 9505 10520
rect 9493 10489 9505 10492
rect 9539 10489 9551 10523
rect 9493 10483 9551 10489
rect 9582 10480 9588 10532
rect 9640 10520 9646 10532
rect 9677 10523 9735 10529
rect 9677 10520 9689 10523
rect 9640 10492 9689 10520
rect 9640 10480 9646 10492
rect 9677 10489 9689 10492
rect 9723 10520 9735 10523
rect 11054 10520 11060 10532
rect 9723 10492 11060 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11333 10523 11391 10529
rect 11333 10489 11345 10523
rect 11379 10520 11391 10523
rect 12544 10520 12572 10551
rect 12618 10548 12624 10600
rect 12676 10588 12682 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 12676 10560 13553 10588
rect 12676 10548 12682 10560
rect 13541 10557 13553 10560
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14384 10588 14412 10764
rect 14918 10616 14924 10668
rect 14976 10616 14982 10668
rect 15102 10588 15108 10600
rect 14231 10560 15108 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 13173 10523 13231 10529
rect 13173 10520 13185 10523
rect 11379 10492 12572 10520
rect 12636 10492 13185 10520
rect 11379 10489 11391 10492
rect 11333 10483 11391 10489
rect 5684 10424 6040 10452
rect 8941 10455 8999 10461
rect 5684 10412 5690 10424
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9030 10452 9036 10464
rect 8987 10424 9036 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11480 10424 11713 10452
rect 11480 10412 11486 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 11882 10412 11888 10464
rect 11940 10412 11946 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12636 10452 12664 10492
rect 13173 10489 13185 10492
rect 13219 10520 13231 10523
rect 14918 10520 14924 10532
rect 13219 10492 14924 10520
rect 13219 10489 13231 10492
rect 13173 10483 13231 10489
rect 14918 10480 14924 10492
rect 14976 10480 14982 10532
rect 12492 10424 12664 10452
rect 12492 10412 12498 10424
rect 12710 10412 12716 10464
rect 12768 10412 12774 10464
rect 12973 10455 13031 10461
rect 12973 10421 12985 10455
rect 13019 10452 13031 10455
rect 13078 10452 13084 10464
rect 13019 10424 13084 10452
rect 13019 10421 13031 10424
rect 12973 10415 13031 10421
rect 13078 10412 13084 10424
rect 13136 10412 13142 10464
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 4614 10208 4620 10260
rect 4672 10248 4678 10260
rect 4709 10251 4767 10257
rect 4709 10248 4721 10251
rect 4672 10220 4721 10248
rect 4672 10208 4678 10220
rect 4709 10217 4721 10220
rect 4755 10217 4767 10251
rect 4709 10211 4767 10217
rect 5258 10208 5264 10260
rect 5316 10208 5322 10260
rect 5718 10208 5724 10260
rect 5776 10248 5782 10260
rect 5813 10251 5871 10257
rect 5813 10248 5825 10251
rect 5776 10220 5825 10248
rect 5776 10208 5782 10220
rect 5813 10217 5825 10220
rect 5859 10217 5871 10251
rect 5813 10211 5871 10217
rect 6181 10251 6239 10257
rect 6181 10217 6193 10251
rect 6227 10248 6239 10251
rect 6454 10248 6460 10260
rect 6227 10220 6460 10248
rect 6227 10217 6239 10220
rect 6181 10211 6239 10217
rect 6454 10208 6460 10220
rect 6512 10248 6518 10260
rect 6914 10248 6920 10260
rect 6512 10220 6920 10248
rect 6512 10208 6518 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10217 7067 10251
rect 7009 10211 7067 10217
rect 8481 10251 8539 10257
rect 8481 10217 8493 10251
rect 8527 10248 8539 10251
rect 8570 10248 8576 10260
rect 8527 10220 8576 10248
rect 8527 10217 8539 10220
rect 8481 10211 8539 10217
rect 4522 10180 4528 10192
rect 4448 10152 4528 10180
rect 4448 10121 4476 10152
rect 4522 10140 4528 10152
rect 4580 10180 4586 10192
rect 5276 10180 5304 10208
rect 6365 10183 6423 10189
rect 6365 10180 6377 10183
rect 4580 10152 6377 10180
rect 4580 10140 4586 10152
rect 6365 10149 6377 10152
rect 6411 10149 6423 10183
rect 7024 10180 7052 10211
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 9398 10248 9404 10260
rect 9048 10220 9404 10248
rect 7346 10183 7404 10189
rect 7346 10180 7358 10183
rect 7024 10152 7358 10180
rect 6365 10143 6423 10149
rect 7346 10149 7358 10152
rect 7392 10149 7404 10183
rect 7346 10143 7404 10149
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 4890 10072 4896 10124
rect 4948 10072 4954 10124
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 5000 10084 5273 10112
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4617 10047 4675 10053
rect 4617 10013 4629 10047
rect 4663 10044 4675 10047
rect 5000 10044 5028 10084
rect 5261 10081 5273 10084
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 5445 10115 5503 10121
rect 5445 10081 5457 10115
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 4663 10016 5028 10044
rect 5077 10047 5135 10053
rect 4663 10013 4675 10016
rect 4617 10007 4675 10013
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5350 10044 5356 10056
rect 5215 10016 5356 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 4264 9908 4292 10007
rect 5092 9976 5120 10007
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5460 10044 5488 10075
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5592 10084 6009 10112
rect 5592 10072 5598 10084
rect 5997 10081 6009 10084
rect 6043 10081 6055 10115
rect 5997 10075 6055 10081
rect 6089 10115 6147 10121
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6546 10112 6552 10124
rect 6135 10084 6552 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 6914 10112 6920 10124
rect 6871 10084 6920 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 8588 10112 8616 10208
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 8588 10084 8769 10112
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 8938 10072 8944 10124
rect 8996 10072 9002 10124
rect 9048 10121 9076 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10192 10220 10609 10248
rect 10192 10208 10198 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 12986 10248 12992 10260
rect 10597 10211 10655 10217
rect 11026 10220 12992 10248
rect 11026 10180 11054 10220
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 9232 10152 11054 10180
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9122 10072 9128 10124
rect 9180 10112 9186 10124
rect 9232 10121 9260 10152
rect 11238 10140 11244 10192
rect 11296 10140 11302 10192
rect 11348 10152 11652 10180
rect 9490 10121 9496 10124
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 9180 10084 9229 10112
rect 9180 10072 9186 10084
rect 9217 10081 9229 10084
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9484 10075 9496 10121
rect 9490 10072 9496 10075
rect 9548 10072 9554 10124
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 11348 10112 11376 10152
rect 11624 10121 11652 10152
rect 11790 10140 11796 10192
rect 11848 10140 11854 10192
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12009 10183 12067 10189
rect 12009 10180 12021 10183
rect 11940 10152 12021 10180
rect 11940 10140 11946 10152
rect 12009 10149 12021 10152
rect 12055 10180 12067 10183
rect 12253 10183 12311 10189
rect 12253 10180 12265 10183
rect 12055 10152 12265 10180
rect 12055 10149 12067 10152
rect 12009 10143 12067 10149
rect 12253 10149 12265 10152
rect 12299 10149 12311 10183
rect 12253 10143 12311 10149
rect 12437 10183 12495 10189
rect 12437 10149 12449 10183
rect 12483 10180 12495 10183
rect 12526 10180 12532 10192
rect 12483 10152 12532 10180
rect 12483 10149 12495 10152
rect 12437 10143 12495 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 12621 10183 12679 10189
rect 12621 10149 12633 10183
rect 12667 10180 12679 10183
rect 12894 10180 12900 10192
rect 12667 10152 12900 10180
rect 12667 10149 12679 10152
rect 12621 10143 12679 10149
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 14645 10183 14703 10189
rect 14645 10149 14657 10183
rect 14691 10180 14703 10183
rect 14918 10180 14924 10192
rect 14691 10152 14924 10180
rect 14691 10149 14703 10152
rect 14645 10143 14703 10149
rect 14918 10140 14924 10152
rect 14976 10140 14982 10192
rect 11204 10084 11376 10112
rect 11425 10115 11483 10121
rect 11204 10072 11210 10084
rect 11425 10081 11437 10115
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 11609 10115 11667 10121
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 12158 10112 12164 10124
rect 11655 10084 12164 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 5460 10016 5764 10044
rect 5626 9976 5632 9988
rect 5092 9948 5632 9976
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5736 9976 5764 10016
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 5868 10016 7113 10044
rect 5868 10004 5874 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 6638 9976 6644 9988
rect 5736 9948 6644 9976
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 11440 9976 11468 10075
rect 12158 10072 12164 10084
rect 12216 10072 12222 10124
rect 12544 10112 12572 10140
rect 12802 10112 12808 10124
rect 12544 10084 12808 10112
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 12986 10072 12992 10124
rect 13044 10072 13050 10124
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10044 11759 10047
rect 11974 10044 11980 10056
rect 11747 10016 11980 10044
rect 11747 10013 11759 10016
rect 11701 10007 11759 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 12768 10016 13277 10044
rect 12768 10004 12774 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 11440 9948 12173 9976
rect 12161 9945 12173 9948
rect 12207 9976 12219 9979
rect 12250 9976 12256 9988
rect 12207 9948 12256 9976
rect 12207 9945 12219 9948
rect 12161 9939 12219 9945
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 8386 9908 8392 9920
rect 4264 9880 8392 9908
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 11514 9868 11520 9920
rect 11572 9868 11578 9920
rect 11977 9911 12035 9917
rect 11977 9877 11989 9911
rect 12023 9908 12035 9911
rect 12526 9908 12532 9920
rect 12023 9880 12532 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 5074 9664 5080 9716
rect 5132 9664 5138 9716
rect 6273 9707 6331 9713
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6546 9704 6552 9716
rect 6319 9676 6552 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6546 9664 6552 9676
rect 6604 9664 6610 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 11609 9707 11667 9713
rect 11609 9704 11621 9707
rect 11572 9676 11621 9704
rect 11572 9664 11578 9676
rect 11609 9673 11621 9676
rect 11655 9673 11667 9707
rect 11609 9667 11667 9673
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 6089 9639 6147 9645
rect 6089 9636 6101 9639
rect 5684 9608 6101 9636
rect 5684 9596 5690 9608
rect 6089 9605 6101 9608
rect 6135 9605 6147 9639
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 6089 9599 6147 9605
rect 7392 9608 8217 9636
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 7392 9577 7420 9608
rect 8205 9605 8217 9608
rect 8251 9636 8263 9639
rect 8478 9636 8484 9648
rect 8251 9608 8484 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 8478 9596 8484 9608
rect 8536 9596 8542 9648
rect 5997 9571 6055 9577
rect 5997 9568 6009 9571
rect 5500 9540 6009 9568
rect 5500 9528 5506 9540
rect 5997 9537 6009 9540
rect 6043 9568 6055 9571
rect 7377 9571 7435 9577
rect 6043 9540 7328 9568
rect 6043 9537 6055 9540
rect 5997 9531 6055 9537
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 5166 9392 5172 9444
rect 5224 9432 5230 9444
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 5224 9404 5273 9432
rect 5224 9392 5230 9404
rect 5261 9401 5273 9404
rect 5307 9432 5319 9435
rect 5442 9432 5448 9444
rect 5307 9404 5448 9432
rect 5307 9401 5319 9404
rect 5261 9395 5319 9401
rect 5442 9392 5448 9404
rect 5500 9392 5506 9444
rect 5552 9432 5580 9463
rect 5626 9460 5632 9512
rect 5684 9460 5690 9512
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9469 7159 9503
rect 7300 9500 7328 9540
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 7708 9540 9229 9568
rect 7708 9528 7714 9540
rect 9217 9537 9229 9540
rect 9263 9537 9275 9571
rect 15010 9568 15016 9580
rect 9217 9531 9275 9537
rect 10980 9540 15016 9568
rect 7466 9500 7472 9512
rect 7300 9472 7472 9500
rect 7101 9463 7159 9469
rect 5718 9432 5724 9444
rect 5552 9404 5724 9432
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 5902 9392 5908 9444
rect 5960 9392 5966 9444
rect 6454 9392 6460 9444
rect 6512 9392 6518 9444
rect 7116 9432 7144 9463
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8938 9500 8944 9512
rect 8067 9472 8944 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 10980 9509 11008 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11333 9503 11391 9509
rect 11333 9469 11345 9503
rect 11379 9500 11391 9503
rect 11422 9500 11428 9512
rect 11379 9472 11428 9500
rect 11379 9469 11391 9472
rect 11333 9463 11391 9469
rect 6748 9404 7144 9432
rect 6748 9376 6776 9404
rect 7558 9392 7564 9444
rect 7616 9432 7622 9444
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7616 9404 7849 9432
rect 7616 9392 7622 9404
rect 7837 9401 7849 9404
rect 7883 9432 7895 9435
rect 10226 9432 10232 9444
rect 7883 9404 10232 9432
rect 7883 9401 7895 9404
rect 7837 9395 7895 9401
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 11348 9432 11376 9463
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 11609 9503 11667 9509
rect 11609 9469 11621 9503
rect 11655 9500 11667 9503
rect 12618 9500 12624 9512
rect 11655 9472 12624 9500
rect 11655 9469 11667 9472
rect 11609 9463 11667 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12802 9460 12808 9512
rect 12860 9460 12866 9512
rect 12989 9503 13047 9509
rect 12989 9469 13001 9503
rect 13035 9500 13047 9503
rect 13078 9500 13084 9512
rect 13035 9472 13084 9500
rect 13035 9469 13047 9472
rect 12989 9463 13047 9469
rect 13078 9460 13084 9472
rect 13136 9500 13142 9512
rect 13541 9503 13599 9509
rect 13541 9500 13553 9503
rect 13136 9472 13553 9500
rect 13136 9460 13142 9472
rect 13541 9469 13553 9472
rect 13587 9469 13599 9503
rect 13541 9463 13599 9469
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9469 13783 9503
rect 13725 9463 13783 9469
rect 13740 9432 13768 9463
rect 13906 9460 13912 9512
rect 13964 9500 13970 9512
rect 14918 9500 14924 9512
rect 13964 9472 14924 9500
rect 13964 9460 13970 9472
rect 14918 9460 14924 9472
rect 14976 9460 14982 9512
rect 13998 9432 14004 9444
rect 11348 9404 12664 9432
rect 13740 9404 14004 9432
rect 12636 9376 12664 9404
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 3878 9324 3884 9376
rect 3936 9364 3942 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 3936 9336 4905 9364
rect 3936 9324 3942 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 5061 9367 5119 9373
rect 5061 9333 5073 9367
rect 5107 9364 5119 9367
rect 5353 9367 5411 9373
rect 5353 9364 5365 9367
rect 5107 9336 5365 9364
rect 5107 9333 5119 9336
rect 5061 9327 5119 9333
rect 5353 9333 5365 9336
rect 5399 9333 5411 9367
rect 5353 9327 5411 9333
rect 6257 9367 6315 9373
rect 6257 9333 6269 9367
rect 6303 9364 6315 9367
rect 6730 9364 6736 9376
rect 6303 9336 6736 9364
rect 6303 9333 6315 9336
rect 6257 9327 6315 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 6822 9324 6828 9376
rect 6880 9324 6886 9376
rect 7098 9324 7104 9376
rect 7156 9364 7162 9376
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 7156 9336 7665 9364
rect 7156 9324 7162 9336
rect 7653 9333 7665 9336
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 7929 9367 7987 9373
rect 7929 9333 7941 9367
rect 7975 9364 7987 9367
rect 9306 9364 9312 9376
rect 7975 9336 9312 9364
rect 7975 9333 7987 9336
rect 7929 9327 7987 9333
rect 9306 9324 9312 9336
rect 9364 9324 9370 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11054 9364 11060 9376
rect 11020 9336 11060 9364
rect 11020 9324 11026 9336
rect 11054 9324 11060 9336
rect 11112 9364 11118 9376
rect 11425 9367 11483 9373
rect 11425 9364 11437 9367
rect 11112 9336 11437 9364
rect 11112 9324 11118 9336
rect 11425 9333 11437 9336
rect 11471 9333 11483 9367
rect 11425 9327 11483 9333
rect 12618 9324 12624 9376
rect 12676 9324 12682 9376
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 4709 9163 4767 9169
rect 4709 9129 4721 9163
rect 4755 9129 4767 9163
rect 4709 9123 4767 9129
rect 4724 9092 4752 9123
rect 5074 9120 5080 9172
rect 5132 9120 5138 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5626 9160 5632 9172
rect 5491 9132 5632 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5626 9120 5632 9132
rect 5684 9160 5690 9172
rect 6546 9160 6552 9172
rect 5684 9132 6552 9160
rect 5684 9120 5690 9132
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7075 9163 7133 9169
rect 7075 9160 7087 9163
rect 6880 9132 7087 9160
rect 6880 9120 6886 9132
rect 7075 9129 7087 9132
rect 7121 9129 7133 9163
rect 7075 9123 7133 9129
rect 8938 9120 8944 9172
rect 8996 9120 9002 9172
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9548 9132 9689 9160
rect 9548 9120 9554 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 10686 9120 10692 9172
rect 10744 9120 10750 9172
rect 13906 9160 13912 9172
rect 13188 9132 13912 9160
rect 5902 9092 5908 9104
rect 4724 9064 5908 9092
rect 3602 9033 3608 9036
rect 3596 8987 3608 9033
rect 3602 8984 3608 8987
rect 3660 8984 3666 9036
rect 5276 9033 5304 9064
rect 5902 9052 5908 9064
rect 5960 9092 5966 9104
rect 6362 9092 6368 9104
rect 5960 9064 6368 9092
rect 5960 9052 5966 9064
rect 6362 9052 6368 9064
rect 6420 9052 6426 9104
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 8754 9092 8760 9104
rect 7340 9064 8760 9092
rect 7340 9052 7346 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 8956 9092 8984 9120
rect 8956 9064 9536 9092
rect 5261 9027 5319 9033
rect 5261 8993 5273 9027
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 5534 8984 5540 9036
rect 5592 8984 5598 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 7006 9024 7012 9036
rect 5776 8996 7012 9024
rect 5776 8984 5782 8996
rect 7006 8984 7012 8996
rect 7064 9024 7070 9036
rect 8846 9024 8852 9036
rect 7064 8996 8852 9024
rect 7064 8984 7070 8996
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 8938 8984 8944 9036
rect 8996 8984 9002 9036
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 9088 8996 9137 9024
rect 9088 8984 9094 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 9214 8984 9220 9036
rect 9272 8984 9278 9036
rect 9309 9027 9367 9033
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 9398 9024 9404 9036
rect 9355 8996 9404 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9508 9033 9536 9064
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 11793 9095 11851 9101
rect 10376 9064 11468 9092
rect 10376 9052 10382 9064
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 10505 9027 10563 9033
rect 10505 8993 10517 9027
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3344 8820 3372 8919
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 7282 8956 7288 8968
rect 5500 8928 7288 8956
rect 5500 8916 5506 8928
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 10520 8956 10548 8987
rect 10686 8984 10692 9036
rect 10744 9024 10750 9036
rect 11440 9033 11468 9064
rect 11793 9061 11805 9095
rect 11839 9092 11851 9095
rect 12802 9092 12808 9104
rect 11839 9064 12808 9092
rect 11839 9061 11851 9064
rect 11793 9055 11851 9061
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 10744 8996 11345 9024
rect 10744 8984 10750 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 8993 11483 9027
rect 11808 9024 11836 9055
rect 12802 9052 12808 9064
rect 12860 9052 12866 9104
rect 11425 8987 11483 8993
rect 11532 8996 11836 9024
rect 7524 8928 10548 8956
rect 7524 8916 7530 8928
rect 6914 8848 6920 8900
rect 6972 8848 6978 8900
rect 10520 8888 10548 8928
rect 10594 8916 10600 8968
rect 10652 8956 10658 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10652 8928 10977 8956
rect 10652 8916 10658 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 10965 8919 11023 8925
rect 11532 8888 11560 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 12529 9027 12587 9033
rect 12529 9024 12541 9027
rect 12492 8996 12541 9024
rect 12492 8984 12498 8996
rect 12529 8993 12541 8996
rect 12575 8993 12587 9027
rect 12529 8987 12587 8993
rect 12710 8984 12716 9036
rect 12768 8984 12774 9036
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 9024 13139 9027
rect 13188 9024 13216 9132
rect 13906 9120 13912 9132
rect 13964 9120 13970 9172
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9061 13323 9095
rect 13265 9055 13323 9061
rect 13127 8996 13216 9024
rect 13280 9024 13308 9055
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13280 8996 13645 9024
rect 13127 8993 13139 8996
rect 13081 8987 13139 8993
rect 13633 8993 13645 8996
rect 13679 8993 13691 9027
rect 13633 8987 13691 8993
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 11655 8928 12817 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8956 12955 8959
rect 12943 8928 13124 8956
rect 12943 8925 12955 8928
rect 12897 8919 12955 8925
rect 13096 8900 13124 8928
rect 13262 8916 13268 8968
rect 13320 8956 13326 8968
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13320 8928 13369 8956
rect 13320 8916 13326 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 10520 8860 11560 8888
rect 13078 8848 13084 8900
rect 13136 8848 13142 8900
rect 3970 8820 3976 8832
rect 3344 8792 3976 8820
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 7101 8823 7159 8829
rect 7101 8789 7113 8823
rect 7147 8820 7159 8823
rect 8570 8820 8576 8832
rect 7147 8792 8576 8820
rect 7147 8789 7159 8792
rect 7101 8783 7159 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 14918 8780 14924 8832
rect 14976 8780 14982 8832
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3697 8619 3755 8625
rect 3697 8616 3709 8619
rect 3660 8588 3709 8616
rect 3660 8576 3666 8588
rect 3697 8585 3709 8588
rect 3743 8585 3755 8619
rect 3697 8579 3755 8585
rect 5353 8619 5411 8625
rect 5353 8585 5365 8619
rect 5399 8616 5411 8619
rect 5626 8616 5632 8628
rect 5399 8588 5632 8616
rect 5399 8585 5411 8588
rect 5353 8579 5411 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 6917 8619 6975 8625
rect 6917 8616 6929 8619
rect 6788 8588 6929 8616
rect 6788 8576 6794 8588
rect 6917 8585 6929 8588
rect 6963 8585 6975 8619
rect 7466 8616 7472 8628
rect 6917 8579 6975 8585
rect 7024 8588 7472 8616
rect 6748 8480 6776 8576
rect 6564 8452 6776 8480
rect 3878 8372 3884 8424
rect 3936 8372 3942 8424
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 6454 8372 6460 8424
rect 6512 8372 6518 8424
rect 6564 8421 6592 8452
rect 6549 8415 6607 8421
rect 6549 8381 6561 8415
rect 6595 8381 6607 8415
rect 6549 8375 6607 8381
rect 6638 8372 6644 8424
rect 6696 8372 6702 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6788 8384 6837 8412
rect 6788 8372 6794 8384
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 7024 8412 7052 8588
rect 7466 8576 7472 8588
rect 7524 8616 7530 8628
rect 8938 8616 8944 8628
rect 7524 8588 8944 8616
rect 7524 8576 7530 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9125 8619 9183 8625
rect 9125 8585 9137 8619
rect 9171 8616 9183 8619
rect 9306 8616 9312 8628
rect 9171 8588 9312 8616
rect 9171 8585 9183 8588
rect 9125 8579 9183 8585
rect 9140 8548 9168 8579
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 12768 8588 13553 8616
rect 12768 8576 12774 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13541 8579 13599 8585
rect 8496 8520 9168 8548
rect 8202 8480 8208 8492
rect 7760 8452 8208 8480
rect 7760 8421 7788 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8386 8440 8392 8492
rect 8444 8440 8450 8492
rect 8496 8489 8524 8520
rect 11422 8508 11428 8560
rect 11480 8508 11486 8560
rect 11701 8551 11759 8557
rect 11701 8517 11713 8551
rect 11747 8548 11759 8551
rect 11885 8551 11943 8557
rect 11885 8548 11897 8551
rect 11747 8520 11897 8548
rect 11747 8517 11759 8520
rect 11701 8511 11759 8517
rect 11885 8517 11897 8520
rect 11931 8517 11943 8551
rect 11885 8511 11943 8517
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 9398 8480 9404 8492
rect 8481 8443 8539 8449
rect 8772 8452 9404 8480
rect 6871 8384 7052 8412
rect 7101 8415 7159 8421
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7745 8415 7803 8421
rect 7745 8412 7757 8415
rect 7331 8384 7757 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7745 8381 7757 8384
rect 7791 8381 7803 8415
rect 7745 8375 7803 8381
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8412 8079 8415
rect 8294 8412 8300 8424
rect 8067 8384 8300 8412
rect 8067 8381 8079 8384
rect 8021 8375 8079 8381
rect 4240 8347 4298 8353
rect 4240 8313 4252 8347
rect 4286 8344 4298 8347
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 4286 8316 6193 8344
rect 4286 8313 4298 8316
rect 4240 8307 4298 8313
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 7116 8288 7144 8375
rect 8294 8372 8300 8384
rect 8352 8412 8358 8424
rect 8496 8412 8524 8443
rect 8352 8384 8524 8412
rect 8352 8372 8358 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8772 8421 8800 8452
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10778 8440 10784 8492
rect 10836 8480 10842 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10836 8452 11529 8480
rect 10836 8440 10842 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 8757 8415 8815 8421
rect 8757 8412 8769 8415
rect 8720 8384 8769 8412
rect 8720 8372 8726 8384
rect 8757 8381 8769 8384
rect 8803 8381 8815 8415
rect 8757 8375 8815 8381
rect 8846 8372 8852 8424
rect 8904 8412 8910 8424
rect 8904 8384 10364 8412
rect 8904 8372 8910 8384
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7837 8347 7895 8353
rect 7837 8344 7849 8347
rect 7616 8316 7849 8344
rect 7616 8304 7622 8316
rect 7837 8313 7849 8316
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 10238 8347 10296 8353
rect 10238 8344 10250 8347
rect 9456 8316 10250 8344
rect 9456 8304 9462 8316
rect 10238 8313 10250 8316
rect 10284 8313 10296 8347
rect 10336 8344 10364 8384
rect 10502 8372 10508 8424
rect 10560 8372 10566 8424
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 11716 8412 11744 8511
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 12529 8483 12587 8489
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 12802 8480 12808 8492
rect 12575 8452 12808 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 11195 8384 11744 8412
rect 11793 8415 11851 8421
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 11793 8381 11805 8415
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 10594 8344 10600 8356
rect 10336 8316 10600 8344
rect 10238 8307 10296 8313
rect 10594 8304 10600 8316
rect 10652 8304 10658 8356
rect 11425 8347 11483 8353
rect 11425 8313 11437 8347
rect 11471 8344 11483 8347
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11471 8316 11529 8344
rect 11471 8313 11483 8316
rect 11425 8307 11483 8313
rect 11517 8313 11529 8316
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 11808 8344 11836 8375
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 13725 8415 13783 8421
rect 13725 8412 13737 8415
rect 12676 8384 13737 8412
rect 12676 8372 12682 8384
rect 13725 8381 13737 8384
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14185 8415 14243 8421
rect 14185 8381 14197 8415
rect 14231 8412 14243 8415
rect 14918 8412 14924 8424
rect 14231 8384 14924 8412
rect 14231 8381 14243 8384
rect 14185 8375 14243 8381
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 13078 8344 13084 8356
rect 11808 8316 13084 8344
rect 5810 8236 5816 8288
rect 5868 8276 5874 8288
rect 7098 8276 7104 8288
rect 5868 8248 7104 8276
rect 5868 8236 5874 8248
rect 7098 8236 7104 8248
rect 7156 8236 7162 8288
rect 8205 8279 8263 8285
rect 8205 8245 8217 8279
rect 8251 8276 8263 8279
rect 8938 8276 8944 8288
rect 8251 8248 8944 8276
rect 8251 8245 8263 8248
rect 8205 8239 8263 8245
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 9030 8236 9036 8288
rect 9088 8236 9094 8288
rect 11146 8236 11152 8288
rect 11204 8276 11210 8288
rect 11241 8279 11299 8285
rect 11241 8276 11253 8279
rect 11204 8248 11253 8276
rect 11204 8236 11210 8248
rect 11241 8245 11253 8248
rect 11287 8276 11299 8279
rect 11808 8276 11836 8316
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 11287 8248 11836 8276
rect 12253 8279 12311 8285
rect 11287 8245 11299 8248
rect 11241 8239 11299 8245
rect 12253 8245 12265 8279
rect 12299 8276 12311 8279
rect 13170 8276 13176 8288
rect 12299 8248 13176 8276
rect 12299 8245 12311 8248
rect 12253 8239 12311 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 7098 8032 7104 8084
rect 7156 8072 7162 8084
rect 7903 8075 7961 8081
rect 7903 8072 7915 8075
rect 7156 8044 7915 8072
rect 7156 8032 7162 8044
rect 7903 8041 7915 8044
rect 7949 8041 7961 8075
rect 7903 8035 7961 8041
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 8497 8075 8555 8081
rect 8497 8072 8509 8075
rect 8260 8044 8509 8072
rect 8260 8032 8266 8044
rect 8497 8041 8509 8044
rect 8543 8041 8555 8075
rect 8497 8035 8555 8041
rect 8662 8032 8668 8084
rect 8720 8032 8726 8084
rect 9398 8032 9404 8084
rect 9456 8032 9462 8084
rect 7650 7964 7656 8016
rect 7708 7964 7714 8016
rect 8113 8007 8171 8013
rect 8113 7973 8125 8007
rect 8159 7973 8171 8007
rect 8113 7967 8171 7973
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 7098 7936 7104 7948
rect 6512 7908 7104 7936
rect 6512 7896 6518 7908
rect 7098 7896 7104 7908
rect 7156 7936 7162 7948
rect 8128 7936 8156 7967
rect 8294 7964 8300 8016
rect 8352 7964 8358 8016
rect 8754 7964 8760 8016
rect 8812 8013 8818 8016
rect 9030 8013 9036 8016
rect 8812 8007 8841 8013
rect 8829 7973 8841 8007
rect 8812 7967 8841 7973
rect 8973 8007 9036 8013
rect 8973 7973 8985 8007
rect 9019 7973 9036 8007
rect 8973 7967 9036 7973
rect 8812 7964 8818 7967
rect 9030 7964 9036 7967
rect 9088 7964 9094 8016
rect 9217 7939 9275 7945
rect 9217 7936 9229 7939
rect 7156 7908 8156 7936
rect 9140 7908 9229 7936
rect 7156 7896 7162 7908
rect 7558 7760 7564 7812
rect 7616 7800 7622 7812
rect 9140 7809 9168 7908
rect 9217 7905 9229 7908
rect 9263 7905 9275 7939
rect 9217 7899 9275 7905
rect 10410 7896 10416 7948
rect 10468 7896 10474 7948
rect 11422 7896 11428 7948
rect 11480 7936 11486 7948
rect 13633 7939 13691 7945
rect 13633 7936 13645 7939
rect 11480 7908 13645 7936
rect 11480 7896 11486 7908
rect 13633 7905 13645 7908
rect 13679 7905 13691 7939
rect 13633 7899 13691 7905
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13262 7868 13268 7880
rect 12952 7840 13268 7868
rect 12952 7828 12958 7840
rect 13262 7828 13268 7840
rect 13320 7868 13326 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 13320 7840 13369 7868
rect 13320 7828 13326 7840
rect 13357 7837 13369 7840
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 9125 7803 9183 7809
rect 7616 7772 8524 7800
rect 7616 7760 7622 7772
rect 8496 7744 8524 7772
rect 9125 7769 9137 7803
rect 9171 7769 9183 7803
rect 9125 7763 9183 7769
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6270 7732 6276 7744
rect 6227 7704 6276 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 6880 7704 7757 7732
rect 6880 7692 6886 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 7745 7695 7803 7701
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8202 7732 8208 7744
rect 7975 7704 8208 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8478 7692 8484 7744
rect 8536 7692 8542 7744
rect 8938 7692 8944 7744
rect 8996 7692 9002 7744
rect 10505 7735 10563 7741
rect 10505 7701 10517 7735
rect 10551 7732 10563 7735
rect 13722 7732 13728 7744
rect 10551 7704 13728 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14734 7692 14740 7744
rect 14792 7692 14798 7744
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 5592 7500 5825 7528
rect 5592 7488 5598 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 6549 7531 6607 7537
rect 6549 7497 6561 7531
rect 6595 7528 6607 7531
rect 6638 7528 6644 7540
rect 6595 7500 6644 7528
rect 6595 7497 6607 7500
rect 6549 7491 6607 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 10686 7528 10692 7540
rect 7208 7500 10692 7528
rect 7208 7404 7236 7500
rect 10686 7488 10692 7500
rect 10744 7528 10750 7540
rect 11238 7528 11244 7540
rect 10744 7500 11244 7528
rect 10744 7488 10750 7500
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 7742 7420 7748 7472
rect 7800 7420 7806 7472
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 12894 7460 12900 7472
rect 10560 7432 12900 7460
rect 10560 7420 10566 7432
rect 12894 7420 12900 7432
rect 12952 7420 12958 7472
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 5776 7364 6745 7392
rect 5776 7352 5782 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6362 7324 6368 7336
rect 5684 7296 6368 7324
rect 5684 7284 5690 7296
rect 6362 7284 6368 7296
rect 6420 7284 6426 7336
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 5997 7259 6055 7265
rect 5997 7256 6009 7259
rect 5868 7228 6009 7256
rect 5868 7216 5874 7228
rect 5997 7225 6009 7228
rect 6043 7225 6055 7259
rect 5997 7219 6055 7225
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6454 7256 6460 7268
rect 6135 7228 6460 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6454 7216 6460 7228
rect 6512 7216 6518 7268
rect 6748 7256 6776 7355
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7650 7352 7656 7404
rect 7708 7392 7714 7404
rect 7708 7364 11652 7392
rect 7708 7352 7714 7364
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 7616 7296 7941 7324
rect 7616 7284 7622 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7324 8079 7327
rect 8202 7324 8208 7336
rect 8067 7296 8208 7324
rect 8067 7293 8079 7296
rect 8021 7287 8079 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 11330 7284 11336 7336
rect 11388 7284 11394 7336
rect 11624 7333 11652 7364
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 14093 7395 14151 7401
rect 14093 7392 14105 7395
rect 12124 7364 14105 7392
rect 12124 7352 12130 7364
rect 14093 7361 14105 7364
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7293 11575 7327
rect 11517 7287 11575 7293
rect 11609 7327 11667 7333
rect 11609 7293 11621 7327
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 6748 7228 7328 7256
rect 5077 7191 5135 7197
rect 5077 7157 5089 7191
rect 5123 7188 5135 7191
rect 5258 7188 5264 7200
rect 5123 7160 5264 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6730 7188 6736 7200
rect 6227 7160 6736 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 7300 7188 7328 7228
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 7745 7259 7803 7265
rect 7745 7256 7757 7259
rect 7432 7228 7757 7256
rect 7432 7216 7438 7228
rect 7745 7225 7757 7228
rect 7791 7225 7803 7259
rect 7745 7219 7803 7225
rect 10962 7216 10968 7268
rect 11020 7256 11026 7268
rect 11532 7256 11560 7287
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 13909 7327 13967 7333
rect 13909 7324 13921 7327
rect 13780 7296 13921 7324
rect 13780 7284 13786 7296
rect 13909 7293 13921 7296
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 11882 7256 11888 7268
rect 11020 7228 11888 7256
rect 11020 7216 11026 7228
rect 11882 7216 11888 7228
rect 11940 7216 11946 7268
rect 11054 7188 11060 7200
rect 7300 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7188 11118 7200
rect 11330 7188 11336 7200
rect 11112 7160 11336 7188
rect 11112 7148 11118 7160
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 12250 7188 12256 7200
rect 11563 7160 12256 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 12250 7148 12256 7160
rect 12308 7148 12314 7200
rect 13538 7148 13544 7200
rect 13596 7148 13602 7200
rect 13998 7148 14004 7200
rect 14056 7148 14062 7200
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 5813 6987 5871 6993
rect 5813 6984 5825 6987
rect 5506 6956 5825 6984
rect 5506 6916 5534 6956
rect 5813 6953 5825 6956
rect 5859 6953 5871 6987
rect 5813 6947 5871 6953
rect 6454 6944 6460 6996
rect 6512 6984 6518 6996
rect 6749 6987 6807 6993
rect 6749 6984 6761 6987
rect 6512 6956 6761 6984
rect 6512 6944 6518 6956
rect 6749 6953 6761 6956
rect 6795 6953 6807 6987
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6749 6947 6807 6953
rect 6840 6956 6929 6984
rect 5460 6888 5534 6916
rect 5460 6860 5488 6888
rect 5718 6876 5724 6928
rect 5776 6916 5782 6928
rect 5776 6888 6040 6916
rect 5776 6876 5782 6888
rect 3688 6851 3746 6857
rect 3688 6817 3700 6851
rect 3734 6848 3746 6851
rect 3734 6820 5028 6848
rect 3734 6817 3746 6820
rect 3688 6811 3746 6817
rect 5000 6789 5028 6820
rect 5258 6808 5264 6860
rect 5316 6808 5322 6860
rect 5353 6851 5411 6857
rect 5353 6817 5365 6851
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5445 6854 5503 6860
rect 5445 6820 5457 6854
rect 5491 6820 5503 6854
rect 5445 6814 5503 6820
rect 5629 6851 5687 6857
rect 5629 6817 5641 6851
rect 5675 6846 5687 6851
rect 5810 6848 5816 6860
rect 5736 6846 5816 6848
rect 5675 6820 5816 6846
rect 5675 6818 5764 6820
rect 5675 6817 5687 6818
rect 5629 6811 5687 6817
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6749 5043 6783
rect 5368 6780 5396 6811
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6012 6857 6040 6888
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 6549 6919 6607 6925
rect 6549 6916 6561 6919
rect 6420 6888 6561 6916
rect 6420 6876 6426 6888
rect 6549 6885 6561 6888
rect 6595 6885 6607 6919
rect 6549 6879 6607 6885
rect 6840 6916 6868 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 9769 6987 9827 6993
rect 9769 6984 9781 6987
rect 8536 6956 9781 6984
rect 8536 6944 8542 6956
rect 9769 6953 9781 6956
rect 9815 6953 9827 6987
rect 9769 6947 9827 6953
rect 10965 6987 11023 6993
rect 10965 6953 10977 6987
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 11425 6987 11483 6993
rect 11425 6953 11437 6987
rect 11471 6984 11483 6987
rect 12066 6984 12072 6996
rect 11471 6956 12072 6984
rect 11471 6953 11483 6956
rect 11425 6947 11483 6953
rect 8202 6916 8208 6928
rect 6840 6888 8208 6916
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6817 6055 6851
rect 5997 6811 6055 6817
rect 6089 6851 6147 6857
rect 6089 6817 6101 6851
rect 6135 6848 6147 6851
rect 6840 6848 6868 6888
rect 6135 6820 6868 6848
rect 6135 6817 6147 6820
rect 6089 6811 6147 6817
rect 5368 6752 5948 6780
rect 4985 6743 5043 6749
rect 3436 6644 3464 6743
rect 5920 6724 5948 6752
rect 5626 6712 5632 6724
rect 4356 6684 5632 6712
rect 4062 6644 4068 6656
rect 3436 6616 4068 6644
rect 4062 6604 4068 6616
rect 4120 6644 4126 6656
rect 4356 6644 4384 6684
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 5902 6672 5908 6724
rect 5960 6672 5966 6724
rect 4120 6616 4384 6644
rect 4801 6647 4859 6653
rect 4120 6604 4126 6616
rect 4801 6613 4813 6647
rect 4847 6644 4859 6647
rect 5488 6644 5494 6656
rect 4847 6616 5494 6644
rect 4847 6613 4859 6616
rect 4801 6607 4859 6613
rect 5488 6604 5494 6616
rect 5546 6604 5552 6656
rect 6012 6644 6040 6811
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7466 6848 7472 6860
rect 6972 6820 7472 6848
rect 6972 6808 6978 6820
rect 7466 6808 7472 6820
rect 7524 6848 7530 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7524 6820 7573 6848
rect 7524 6808 7530 6820
rect 7561 6817 7573 6820
rect 7607 6817 7619 6851
rect 7561 6811 7619 6817
rect 7742 6808 7748 6860
rect 7800 6808 7806 6860
rect 7944 6857 7972 6888
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 8297 6919 8355 6925
rect 8297 6885 8309 6919
rect 8343 6916 8355 6919
rect 8634 6919 8692 6925
rect 8634 6916 8646 6919
rect 8343 6888 8646 6916
rect 8343 6885 8355 6888
rect 8297 6879 8355 6885
rect 8634 6885 8646 6888
rect 8680 6885 8692 6919
rect 8634 6879 8692 6885
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8478 6848 8484 6860
rect 8159 6820 8484 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6817 10195 6851
rect 10137 6811 10195 6817
rect 10321 6851 10379 6857
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 10980 6848 11008 6947
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13170 6984 13176 6996
rect 13004 6956 13176 6984
rect 11882 6876 11888 6928
rect 11940 6916 11946 6928
rect 11940 6888 12756 6916
rect 11940 6876 11946 6888
rect 10367 6820 11008 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6546 6780 6552 6792
rect 6503 6752 6552 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6546 6740 6552 6752
rect 6604 6780 6610 6792
rect 7190 6780 7196 6792
rect 6604 6752 7196 6780
rect 6604 6740 6610 6752
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7708 6752 7849 6780
rect 7708 6740 7714 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8386 6740 8392 6792
rect 8444 6740 8450 6792
rect 6270 6672 6276 6724
rect 6328 6712 6334 6724
rect 8404 6712 8432 6740
rect 6328 6684 8432 6712
rect 10152 6712 10180 6811
rect 11330 6808 11336 6860
rect 11388 6848 11394 6860
rect 12161 6851 12219 6857
rect 11388 6820 12112 6848
rect 11388 6808 11394 6820
rect 12084 6792 12112 6820
rect 12161 6817 12173 6851
rect 12207 6848 12219 6851
rect 12434 6848 12440 6860
rect 12207 6820 12440 6848
rect 12207 6817 12219 6820
rect 12161 6811 12219 6817
rect 12434 6808 12440 6820
rect 12492 6848 12498 6860
rect 12728 6857 12756 6888
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12492 6820 12541 6848
rect 12492 6808 12498 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12713 6851 12771 6857
rect 12713 6817 12725 6851
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 12894 6808 12900 6860
rect 12952 6808 12958 6860
rect 13004 6857 13032 6956
rect 13170 6944 13176 6956
rect 13228 6984 13234 6996
rect 14734 6984 14740 6996
rect 13228 6956 14740 6984
rect 13228 6944 13234 6956
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 13538 6876 13544 6928
rect 13596 6876 13602 6928
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6817 13047 6851
rect 12989 6811 13047 6817
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 13136 6820 13461 6848
rect 13136 6808 13142 6820
rect 13449 6817 13461 6820
rect 13495 6848 13507 6851
rect 13722 6848 13728 6860
rect 13495 6820 13728 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 11054 6740 11060 6792
rect 11112 6780 11118 6792
rect 11517 6783 11575 6789
rect 11517 6780 11529 6783
rect 11112 6752 11529 6780
rect 11112 6740 11118 6752
rect 11517 6749 11529 6752
rect 11563 6749 11575 6783
rect 11517 6743 11575 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 10152 6684 11054 6712
rect 6328 6672 6334 6684
rect 6454 6644 6460 6656
rect 6012 6616 6460 6644
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 6730 6604 6736 6656
rect 6788 6604 6794 6656
rect 10318 6604 10324 6656
rect 10376 6604 10382 6656
rect 11026 6644 11054 6684
rect 11992 6644 12020 6743
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12250 6740 12256 6792
rect 12308 6740 12314 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 12400 6752 13185 6780
rect 12400 6740 12406 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13173 6743 13231 6749
rect 12710 6672 12716 6724
rect 12768 6712 12774 6724
rect 13265 6715 13323 6721
rect 13265 6712 13277 6715
rect 12768 6684 13277 6712
rect 12768 6672 12774 6684
rect 13265 6681 13277 6684
rect 13311 6681 13323 6715
rect 13265 6675 13323 6681
rect 12158 6644 12164 6656
rect 11026 6616 12164 6644
rect 12158 6604 12164 6616
rect 12216 6644 12222 6656
rect 12342 6644 12348 6656
rect 12216 6616 12348 6644
rect 12216 6604 12222 6616
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12618 6644 12624 6656
rect 12483 6616 12624 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 13078 6604 13084 6656
rect 13136 6604 13142 6656
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 6270 6440 6276 6452
rect 5684 6412 6276 6440
rect 5684 6400 5690 6412
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6440 7343 6443
rect 7374 6440 7380 6452
rect 7331 6412 7380 6440
rect 7331 6409 7343 6412
rect 7285 6403 7343 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7653 6443 7711 6449
rect 7653 6409 7665 6443
rect 7699 6440 7711 6443
rect 7742 6440 7748 6452
rect 7699 6412 7748 6440
rect 7699 6409 7711 6412
rect 7653 6403 7711 6409
rect 7742 6400 7748 6412
rect 7800 6400 7806 6452
rect 12710 6400 12716 6452
rect 12768 6400 12774 6452
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 12952 6412 13185 6440
rect 12952 6400 12958 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 13998 6440 14004 6452
rect 13403 6412 14004 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 4801 6375 4859 6381
rect 4801 6341 4813 6375
rect 4847 6372 4859 6375
rect 5994 6372 6000 6384
rect 4847 6344 6000 6372
rect 4847 6341 4859 6344
rect 4801 6335 4859 6341
rect 5994 6332 6000 6344
rect 6052 6372 6058 6384
rect 6730 6372 6736 6384
rect 6052 6344 6736 6372
rect 6052 6332 6058 6344
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 6454 6304 6460 6316
rect 5675 6276 6460 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6564 6313 6592 6344
rect 6730 6332 6736 6344
rect 6788 6332 6794 6384
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6638 6264 6644 6316
rect 6696 6304 6702 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 6696 6276 8033 6304
rect 6696 6264 6702 6276
rect 8021 6273 8033 6276
rect 8067 6304 8079 6307
rect 8294 6304 8300 6316
rect 8067 6276 8300 6304
rect 8067 6273 8079 6276
rect 8021 6267 8079 6273
rect 8294 6264 8300 6276
rect 8352 6304 8358 6316
rect 9122 6304 9128 6316
rect 8352 6276 9128 6304
rect 8352 6264 8358 6276
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3970 6236 3976 6248
rect 3467 6208 3976 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3970 6196 3976 6208
rect 4028 6196 4034 6248
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 6181 6239 6239 6245
rect 6181 6236 6193 6239
rect 5776 6208 6193 6236
rect 5776 6196 5782 6208
rect 6181 6205 6193 6208
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 6362 6196 6368 6248
rect 6420 6196 6426 6248
rect 7098 6196 7104 6248
rect 7156 6196 7162 6248
rect 7558 6196 7564 6248
rect 7616 6236 7622 6248
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 7616 6208 7849 6236
rect 7616 6196 7622 6208
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 9456 6208 9781 6236
rect 9456 6196 9462 6208
rect 9769 6205 9781 6208
rect 9815 6236 9827 6239
rect 10502 6236 10508 6248
rect 9815 6208 10508 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 10502 6196 10508 6208
rect 10560 6196 10566 6248
rect 12434 6196 12440 6248
rect 12492 6196 12498 6248
rect 12713 6239 12771 6245
rect 12713 6205 12725 6239
rect 12759 6236 12771 6239
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 12759 6208 13829 6236
rect 12759 6205 12771 6208
rect 12713 6199 12771 6205
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 14461 6239 14519 6245
rect 14461 6205 14473 6239
rect 14507 6236 14519 6239
rect 14918 6236 14924 6248
rect 14507 6208 14924 6236
rect 14507 6205 14519 6208
rect 14461 6199 14519 6205
rect 3688 6171 3746 6177
rect 3688 6137 3700 6171
rect 3734 6168 3746 6171
rect 4890 6168 4896 6180
rect 3734 6140 4896 6168
rect 3734 6137 3746 6140
rect 3688 6131 3746 6137
rect 4890 6128 4896 6140
rect 4948 6128 4954 6180
rect 5994 6128 6000 6180
rect 6052 6128 6058 6180
rect 6089 6171 6147 6177
rect 6089 6137 6101 6171
rect 6135 6168 6147 6171
rect 6546 6168 6552 6180
rect 6135 6140 6552 6168
rect 6135 6137 6147 6140
rect 6089 6131 6147 6137
rect 6546 6128 6552 6140
rect 6604 6128 6610 6180
rect 10036 6171 10094 6177
rect 10036 6137 10048 6171
rect 10082 6168 10094 6171
rect 10318 6168 10324 6180
rect 10082 6140 10324 6168
rect 10082 6137 10094 6140
rect 10036 6131 10094 6137
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 12989 6171 13047 6177
rect 12989 6137 13001 6171
rect 13035 6168 13047 6171
rect 14476 6168 14504 6199
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 13035 6140 14504 6168
rect 13035 6137 13047 6140
rect 12989 6131 13047 6137
rect 5350 6060 5356 6112
rect 5408 6100 5414 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 5408 6072 5457 6100
rect 5408 6060 5414 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 11112 6072 11161 6100
rect 11112 6060 11118 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11149 6063 11207 6069
rect 12066 6060 12072 6112
rect 12124 6100 12130 6112
rect 12434 6100 12440 6112
rect 12124 6072 12440 6100
rect 12124 6060 12130 6072
rect 12434 6060 12440 6072
rect 12492 6100 12498 6112
rect 12529 6103 12587 6109
rect 12529 6100 12541 6103
rect 12492 6072 12541 6100
rect 12492 6060 12498 6072
rect 12529 6069 12541 6072
rect 12575 6069 12587 6103
rect 12529 6063 12587 6069
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 13170 6100 13176 6112
rect 13228 6109 13234 6112
rect 13228 6103 13247 6109
rect 12860 6072 13176 6100
rect 12860 6060 12866 6072
rect 13170 6060 13176 6072
rect 13235 6100 13247 6103
rect 13814 6100 13820 6112
rect 13235 6072 13820 6100
rect 13235 6069 13247 6072
rect 13228 6063 13247 6069
rect 13228 6060 13234 6063
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 8938 5896 8944 5908
rect 7852 5868 8944 5896
rect 6638 5828 6644 5840
rect 6380 5800 6644 5828
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5994 5760 6000 5772
rect 5675 5732 6000 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 6270 5720 6276 5772
rect 6328 5760 6334 5772
rect 6380 5769 6408 5800
rect 6638 5788 6644 5800
rect 6696 5788 6702 5840
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 7561 5831 7619 5837
rect 7561 5828 7573 5831
rect 7432 5800 7573 5828
rect 7432 5788 7438 5800
rect 7561 5797 7573 5800
rect 7607 5797 7619 5831
rect 7561 5791 7619 5797
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 6328 5732 6377 5760
rect 6328 5720 6334 5732
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6730 5760 6736 5772
rect 6503 5732 6736 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6730 5720 6736 5732
rect 6788 5760 6794 5772
rect 7742 5760 7748 5772
rect 6788 5732 7748 5760
rect 6788 5720 6794 5732
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 7852 5769 7880 5868
rect 8938 5856 8944 5868
rect 8996 5896 9002 5908
rect 9585 5899 9643 5905
rect 9585 5896 9597 5899
rect 8996 5868 9597 5896
rect 8996 5856 9002 5868
rect 9585 5865 9597 5868
rect 9631 5865 9643 5899
rect 10778 5896 10784 5908
rect 9585 5859 9643 5865
rect 9692 5868 10784 5896
rect 8662 5837 8668 5840
rect 8649 5831 8668 5837
rect 8649 5797 8661 5831
rect 8649 5791 8668 5797
rect 8662 5788 8668 5791
rect 8720 5788 8726 5840
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 8849 5831 8907 5837
rect 8849 5828 8861 5831
rect 8812 5800 8861 5828
rect 8812 5788 8818 5800
rect 8849 5797 8861 5800
rect 8895 5828 8907 5831
rect 9692 5828 9720 5868
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11480 5868 11897 5896
rect 11480 5856 11486 5868
rect 11885 5865 11897 5868
rect 11931 5896 11943 5899
rect 11974 5896 11980 5908
rect 11931 5868 11980 5896
rect 11931 5865 11943 5868
rect 11885 5859 11943 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 8895 5800 9720 5828
rect 9861 5831 9919 5837
rect 8895 5797 8907 5800
rect 8849 5791 8907 5797
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 10318 5828 10324 5840
rect 9907 5800 10324 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 10318 5788 10324 5800
rect 10376 5788 10382 5840
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5729 7895 5763
rect 7837 5723 7895 5729
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5760 8079 5763
rect 9769 5763 9827 5769
rect 8067 5732 8524 5760
rect 8067 5729 8079 5732
rect 8021 5723 8079 5729
rect 5718 5584 5724 5636
rect 5776 5624 5782 5636
rect 6822 5624 6828 5636
rect 5776 5596 6828 5624
rect 5776 5584 5782 5596
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 8496 5633 8524 5732
rect 9769 5729 9781 5763
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 9953 5763 10011 5769
rect 9953 5729 9965 5763
rect 9999 5760 10011 5763
rect 10042 5760 10048 5772
rect 9999 5732 10048 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 9784 5692 9812 5723
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10796 5760 10824 5856
rect 11701 5763 11759 5769
rect 11701 5760 11713 5763
rect 10796 5732 11713 5760
rect 11701 5729 11713 5732
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 12713 5763 12771 5769
rect 12713 5760 12725 5763
rect 12676 5732 12725 5760
rect 12676 5720 12682 5732
rect 12713 5729 12725 5732
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 12986 5720 12992 5772
rect 13044 5720 13050 5772
rect 13170 5720 13176 5772
rect 13228 5720 13234 5772
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 13357 5763 13415 5769
rect 13357 5760 13369 5763
rect 13320 5732 13369 5760
rect 13320 5720 13326 5732
rect 13357 5729 13369 5732
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 9784 5664 10272 5692
rect 8481 5627 8539 5633
rect 8481 5593 8493 5627
rect 8527 5593 8539 5627
rect 8481 5587 8539 5593
rect 10134 5584 10140 5636
rect 10192 5584 10198 5636
rect 10244 5568 10272 5664
rect 13078 5652 13084 5704
rect 13136 5692 13142 5704
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 13136 5664 13645 5692
rect 13136 5652 13142 5664
rect 13633 5661 13645 5664
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5166 5556 5172 5568
rect 5031 5528 5172 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 6641 5559 6699 5565
rect 6641 5525 6653 5559
rect 6687 5556 6699 5559
rect 6914 5556 6920 5568
rect 6687 5528 6920 5556
rect 6687 5525 6699 5528
rect 6641 5519 6699 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 7064 5528 7573 5556
rect 7064 5516 7070 5528
rect 7561 5525 7573 5528
rect 7607 5525 7619 5559
rect 7561 5519 7619 5525
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8294 5556 8300 5568
rect 8251 5528 8300 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8665 5559 8723 5565
rect 8665 5525 8677 5559
rect 8711 5556 8723 5559
rect 9306 5556 9312 5568
rect 8711 5528 9312 5556
rect 8711 5525 8723 5528
rect 8665 5519 8723 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 10226 5516 10232 5568
rect 10284 5556 10290 5568
rect 11054 5556 11060 5568
rect 10284 5528 11060 5556
rect 10284 5516 10290 5528
rect 11054 5516 11060 5528
rect 11112 5556 11118 5568
rect 11790 5556 11796 5568
rect 11112 5528 11796 5556
rect 11112 5516 11118 5528
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 12529 5559 12587 5565
rect 12529 5525 12541 5559
rect 12575 5556 12587 5559
rect 13078 5556 13084 5568
rect 12575 5528 13084 5556
rect 12575 5525 12587 5528
rect 12529 5519 12587 5525
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 14918 5516 14924 5568
rect 14976 5556 14982 5568
rect 15654 5556 15660 5568
rect 14976 5528 15660 5556
rect 14976 5516 14982 5528
rect 15654 5516 15660 5528
rect 15712 5516 15718 5568
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 4890 5312 4896 5364
rect 4948 5312 4954 5364
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 10318 5352 10324 5364
rect 10091 5324 10324 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 11296 5324 12756 5352
rect 11296 5312 11302 5324
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 7098 5284 7104 5296
rect 5868 5256 7104 5284
rect 5868 5244 5874 5256
rect 7098 5244 7104 5256
rect 7156 5284 7162 5296
rect 8202 5284 8208 5296
rect 7156 5256 8208 5284
rect 7156 5244 7162 5256
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 9769 5287 9827 5293
rect 9769 5253 9781 5287
rect 9815 5284 9827 5287
rect 10134 5284 10140 5296
rect 9815 5256 10140 5284
rect 9815 5253 9827 5256
rect 9769 5247 9827 5253
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 10229 5287 10287 5293
rect 10229 5253 10241 5287
rect 10275 5253 10287 5287
rect 12529 5287 12587 5293
rect 12529 5284 12541 5287
rect 10229 5247 10287 5253
rect 11716 5256 12541 5284
rect 5276 5188 5948 5216
rect 5166 5108 5172 5160
rect 5224 5108 5230 5160
rect 5276 5157 5304 5188
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5350 5108 5356 5160
rect 5408 5108 5414 5160
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 5718 5148 5724 5160
rect 5583 5120 5724 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5810 5108 5816 5160
rect 5868 5108 5874 5160
rect 5920 5157 5948 5188
rect 6270 5176 6276 5228
rect 6328 5176 6334 5228
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7742 5176 7748 5228
rect 7800 5216 7806 5228
rect 8113 5219 8171 5225
rect 8113 5216 8125 5219
rect 7800 5188 8125 5216
rect 7800 5176 7806 5188
rect 8113 5185 8125 5188
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 10042 5176 10048 5228
rect 10100 5176 10106 5228
rect 10244 5216 10272 5247
rect 10244 5188 10640 5216
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5148 5963 5151
rect 6362 5148 6368 5160
rect 5951 5120 6368 5148
rect 5951 5117 5963 5120
rect 5905 5111 5963 5117
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 6822 5148 6828 5160
rect 6779 5120 6828 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 6914 5108 6920 5160
rect 6972 5108 6978 5160
rect 7098 5108 7104 5160
rect 7156 5157 7162 5160
rect 7156 5151 7205 5157
rect 7156 5117 7159 5151
rect 7193 5117 7205 5151
rect 7156 5111 7205 5117
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5148 7343 5151
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7331 5120 7573 5148
rect 7331 5117 7343 5120
rect 7285 5111 7343 5117
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 7561 5111 7619 5117
rect 7156 5108 7162 5111
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8645 5151 8703 5157
rect 8645 5148 8657 5151
rect 8352 5120 8657 5148
rect 8352 5108 8358 5120
rect 8645 5117 8657 5120
rect 8691 5117 8703 5151
rect 10060 5148 10088 5176
rect 8645 5111 8703 5117
rect 9876 5120 10364 5148
rect 5994 5040 6000 5092
rect 6052 5080 6058 5092
rect 6181 5083 6239 5089
rect 6181 5080 6193 5083
rect 6052 5052 6193 5080
rect 6052 5040 6058 5052
rect 6181 5049 6193 5052
rect 6227 5049 6239 5083
rect 6181 5043 6239 5049
rect 9766 5040 9772 5092
rect 9824 5080 9830 5092
rect 9876 5089 9904 5120
rect 9861 5083 9919 5089
rect 9861 5080 9873 5083
rect 9824 5052 9873 5080
rect 9824 5040 9830 5052
rect 9861 5049 9873 5052
rect 9907 5049 9919 5083
rect 9861 5043 9919 5049
rect 10077 5083 10135 5089
rect 10077 5049 10089 5083
rect 10123 5080 10135 5083
rect 10226 5080 10232 5092
rect 10123 5052 10232 5080
rect 10123 5049 10135 5052
rect 10077 5043 10135 5049
rect 10226 5040 10232 5052
rect 10284 5040 10290 5092
rect 10336 5080 10364 5120
rect 10502 5108 10508 5160
rect 10560 5108 10566 5160
rect 10612 5157 10640 5188
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 11716 5225 11744 5256
rect 12529 5253 12541 5256
rect 12575 5253 12587 5287
rect 12529 5247 12587 5253
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 12728 5225 12756 5324
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 13044 5324 13185 5352
rect 13044 5312 13050 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 12894 5244 12900 5296
rect 12952 5284 12958 5296
rect 12952 5256 14596 5284
rect 12952 5244 12958 5256
rect 12713 5219 12771 5225
rect 11848 5188 12296 5216
rect 11848 5176 11854 5188
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 11422 5108 11428 5160
rect 11480 5108 11486 5160
rect 12268 5157 12296 5188
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 13170 5176 13176 5228
rect 13228 5216 13234 5228
rect 14568 5225 14596 5256
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13228 5188 14013 5216
rect 13228 5176 13234 5188
rect 14001 5185 14013 5188
rect 14047 5185 14059 5219
rect 14001 5179 14059 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 14642 5216 14648 5228
rect 14599 5188 14648 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5117 11667 5151
rect 11609 5111 11667 5117
rect 11988 5151 12046 5157
rect 11988 5117 12000 5151
rect 12034 5148 12046 5151
rect 12253 5151 12311 5157
rect 12034 5120 12112 5148
rect 12034 5117 12046 5120
rect 11988 5111 12046 5117
rect 10873 5083 10931 5089
rect 10336 5052 10548 5080
rect 10520 5024 10548 5052
rect 10873 5049 10885 5083
rect 10919 5049 10931 5083
rect 11624 5080 11652 5111
rect 11882 5080 11888 5092
rect 11624 5052 11888 5080
rect 10873 5043 10931 5049
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 7466 4972 7472 5024
rect 7524 4972 7530 5024
rect 10318 4972 10324 5024
rect 10376 4972 10382 5024
rect 10502 4972 10508 5024
rect 10560 5012 10566 5024
rect 10888 5012 10916 5043
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12084 5080 12112 5120
rect 12253 5117 12265 5151
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12492 5120 13001 5148
rect 12492 5108 12498 5120
rect 12989 5117 13001 5120
rect 13035 5117 13047 5151
rect 12989 5111 13047 5117
rect 12345 5083 12403 5089
rect 12345 5080 12357 5083
rect 12084 5052 12357 5080
rect 12084 5024 12112 5052
rect 12345 5049 12357 5052
rect 12391 5049 12403 5083
rect 12345 5043 12403 5049
rect 12529 5083 12587 5089
rect 12529 5049 12541 5083
rect 12575 5080 12587 5083
rect 13722 5080 13728 5092
rect 12575 5052 13728 5080
rect 12575 5049 12587 5052
rect 12529 5043 12587 5049
rect 13722 5040 13728 5052
rect 13780 5040 13786 5092
rect 10560 4984 10916 5012
rect 10560 4972 10566 4984
rect 12066 4972 12072 5024
rect 12124 4972 12130 5024
rect 12158 4972 12164 5024
rect 12216 4972 12222 5024
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5718 4808 5724 4820
rect 5491 4780 5724 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5718 4768 5724 4780
rect 5776 4808 5782 4820
rect 5994 4808 6000 4820
rect 5776 4780 6000 4808
rect 5776 4768 5782 4780
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6270 4808 6276 4820
rect 6227 4780 6276 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6270 4768 6276 4780
rect 6328 4808 6334 4820
rect 6730 4808 6736 4820
rect 6328 4780 6736 4808
rect 6328 4768 6334 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 8662 4768 8668 4820
rect 8720 4768 8726 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9364 4780 9413 4808
rect 9364 4768 9370 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10410 4808 10416 4820
rect 9732 4780 10416 4808
rect 9732 4768 9738 4780
rect 10410 4768 10416 4780
rect 10468 4808 10474 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 10468 4780 10609 4808
rect 10468 4768 10474 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 11882 4808 11888 4820
rect 11747 4780 11888 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 7466 4700 7472 4752
rect 7524 4740 7530 4752
rect 7846 4743 7904 4749
rect 7846 4740 7858 4743
rect 7524 4712 7858 4740
rect 7524 4700 7530 4712
rect 7846 4709 7858 4712
rect 7892 4709 7904 4743
rect 10612 4740 10640 4771
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 14642 4768 14648 4820
rect 14700 4768 14706 4820
rect 7846 4703 7904 4709
rect 7944 4712 8984 4740
rect 10612 4712 11560 4740
rect 3970 4632 3976 4684
rect 4028 4672 4034 4684
rect 4338 4681 4344 4684
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 4028 4644 4077 4672
rect 4028 4632 4034 4644
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 4332 4635 4344 4681
rect 4338 4632 4344 4635
rect 4396 4632 4402 4684
rect 5994 4632 6000 4684
rect 6052 4632 6058 4684
rect 6273 4675 6331 4681
rect 6273 4641 6285 4675
rect 6319 4672 6331 4675
rect 6454 4672 6460 4684
rect 6319 4644 6460 4672
rect 6319 4641 6331 4644
rect 6273 4635 6331 4641
rect 6454 4632 6460 4644
rect 6512 4672 6518 4684
rect 7098 4672 7104 4684
rect 6512 4644 7104 4672
rect 6512 4632 6518 4644
rect 7098 4632 7104 4644
rect 7156 4672 7162 4684
rect 7944 4672 7972 4712
rect 8956 4684 8984 4712
rect 7156 4644 7972 4672
rect 8113 4675 8171 4681
rect 7156 4632 7162 4644
rect 8113 4641 8125 4675
rect 8159 4672 8171 4675
rect 8386 4672 8392 4684
rect 8159 4644 8392 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 8938 4632 8944 4684
rect 8996 4632 9002 4684
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 9180 4644 9321 4672
rect 9180 4632 9186 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 9309 4635 9367 4641
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 10226 4672 10232 4684
rect 9631 4644 10232 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 10502 4672 10508 4684
rect 10459 4644 10508 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 11054 4672 11060 4684
rect 10735 4644 11060 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11532 4681 11560 4712
rect 12158 4700 12164 4752
rect 12216 4740 12222 4752
rect 12906 4743 12964 4749
rect 12906 4740 12918 4743
rect 12216 4712 12918 4740
rect 12216 4700 12222 4712
rect 12906 4709 12918 4712
rect 12952 4709 12964 4743
rect 12906 4703 12964 4709
rect 13078 4700 13084 4752
rect 13136 4740 13142 4752
rect 13136 4712 13400 4740
rect 13136 4700 13142 4712
rect 11333 4675 11391 4681
rect 11333 4672 11345 4675
rect 11296 4644 11345 4672
rect 11296 4632 11302 4644
rect 11333 4641 11345 4644
rect 11379 4641 11391 4675
rect 11333 4635 11391 4641
rect 11517 4675 11575 4681
rect 11517 4641 11529 4675
rect 11563 4672 11575 4675
rect 13173 4675 13231 4681
rect 11563 4644 11836 4672
rect 11563 4641 11575 4644
rect 11517 4635 11575 4641
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 8849 4607 8907 4613
rect 8849 4604 8861 4607
rect 8260 4576 8861 4604
rect 8260 4564 8266 4576
rect 8849 4573 8861 4576
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9232 4536 9260 4567
rect 9674 4564 9680 4616
rect 9732 4564 9738 4616
rect 9766 4564 9772 4616
rect 9824 4564 9830 4616
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 10134 4604 10140 4616
rect 9907 4576 10140 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 9876 4536 9904 4567
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 11808 4545 11836 4644
rect 13173 4641 13185 4675
rect 13219 4672 13231 4675
rect 13262 4672 13268 4684
rect 13219 4644 13268 4672
rect 13219 4641 13231 4644
rect 13173 4635 13231 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13372 4672 13400 4712
rect 13541 4675 13599 4681
rect 13541 4672 13553 4675
rect 13372 4644 13553 4672
rect 13541 4641 13553 4644
rect 13587 4641 13599 4675
rect 13541 4635 13599 4641
rect 9232 4508 9904 4536
rect 11793 4539 11851 4545
rect 11793 4505 11805 4539
rect 11839 4536 11851 4539
rect 12066 4536 12072 4548
rect 11839 4508 12072 4536
rect 11839 4505 11851 4508
rect 11793 4499 11851 4505
rect 12066 4496 12072 4508
rect 12124 4496 12130 4548
rect 5810 4428 5816 4480
rect 5868 4428 5874 4480
rect 10226 4428 10232 4480
rect 10284 4428 10290 4480
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 4396 4236 4445 4264
rect 4396 4224 4402 4236
rect 4433 4233 4445 4236
rect 4479 4233 4491 4267
rect 4433 4227 4491 4233
rect 5169 4267 5227 4273
rect 5169 4233 5181 4267
rect 5215 4264 5227 4267
rect 5810 4264 5816 4276
rect 5215 4236 5816 4264
rect 5215 4233 5227 4236
rect 5169 4227 5227 4233
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 6270 4264 6276 4276
rect 6135 4236 6276 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 10226 4224 10232 4276
rect 10284 4224 10290 4276
rect 4617 4063 4675 4069
rect 4617 4029 4629 4063
rect 4663 4060 4675 4063
rect 8754 4060 8760 4072
rect 4663 4032 5028 4060
rect 4663 4029 4675 4032
rect 4617 4023 4675 4029
rect 5000 3933 5028 4032
rect 5368 4032 8760 4060
rect 5368 4001 5396 4032
rect 8754 4020 8760 4032
rect 8812 4060 8818 4072
rect 8812 4032 10088 4060
rect 8812 4020 8818 4032
rect 5353 3995 5411 4001
rect 5353 3961 5365 3995
rect 5399 3961 5411 3995
rect 5353 3955 5411 3961
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 5905 3995 5963 4001
rect 5905 3992 5917 3995
rect 5776 3964 5917 3992
rect 5776 3952 5782 3964
rect 5905 3961 5917 3964
rect 5951 3961 5963 3995
rect 5905 3955 5963 3961
rect 6121 3995 6179 4001
rect 6121 3961 6133 3995
rect 6167 3992 6179 3995
rect 6454 3992 6460 4004
rect 6167 3964 6460 3992
rect 6167 3961 6179 3964
rect 6121 3955 6179 3961
rect 6454 3952 6460 3964
rect 6512 3952 6518 4004
rect 10060 4001 10088 4032
rect 10318 4001 10324 4004
rect 10045 3995 10103 4001
rect 10045 3961 10057 3995
rect 10091 3961 10103 3995
rect 10045 3955 10103 3961
rect 10261 3995 10324 4001
rect 10261 3961 10273 3995
rect 10307 3961 10324 3995
rect 10261 3955 10324 3961
rect 10318 3952 10324 3955
rect 10376 3952 10382 4004
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3893 5043 3927
rect 4985 3887 5043 3893
rect 5153 3927 5211 3933
rect 5153 3893 5165 3927
rect 5199 3924 5211 3927
rect 5626 3924 5632 3936
rect 5199 3896 5632 3924
rect 5199 3893 5211 3896
rect 5153 3887 5211 3893
rect 5626 3884 5632 3896
rect 5684 3884 5690 3936
rect 6273 3927 6331 3933
rect 6273 3893 6285 3927
rect 6319 3924 6331 3927
rect 6362 3924 6368 3936
rect 6319 3896 6368 3924
rect 6319 3893 6331 3896
rect 6273 3887 6331 3893
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 10410 3884 10416 3936
rect 10468 3884 10474 3936
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 10502 3680 10508 3732
rect 10560 3720 10566 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10560 3692 10793 3720
rect 10560 3680 10566 3692
rect 10781 3689 10793 3692
rect 10827 3689 10839 3723
rect 10781 3683 10839 3689
rect 9398 3544 9404 3596
rect 9456 3544 9462 3596
rect 9668 3587 9726 3593
rect 9668 3553 9680 3587
rect 9714 3584 9726 3587
rect 10042 3584 10048 3596
rect 9714 3556 10048 3584
rect 9714 3553 9726 3556
rect 9668 3547 9726 3553
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 10042 3136 10048 3188
rect 10100 3136 10106 3188
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 10410 2972 10416 2984
rect 10275 2944 10416 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
<< via1 >>
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 5080 15036 5132 15088
rect 940 15011 992 15020
rect 940 14977 949 15011
rect 949 14977 983 15011
rect 983 14977 992 15011
rect 940 14968 992 14977
rect 4436 14968 4488 15020
rect 2136 14900 2188 14952
rect 3516 14943 3568 14952
rect 3516 14909 3525 14943
rect 3525 14909 3559 14943
rect 3559 14909 3568 14943
rect 3516 14900 3568 14909
rect 4620 14900 4672 14952
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 5816 14900 5868 14952
rect 7288 14900 7340 14952
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 9220 14943 9272 14952
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 10048 14900 10100 14952
rect 11152 14900 11204 14952
rect 12440 14900 12492 14952
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 13728 14900 13780 14952
rect 3608 14764 3660 14816
rect 4712 14764 4764 14816
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 6368 14764 6420 14816
rect 6920 14764 6972 14816
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 8944 14764 8996 14816
rect 10416 14764 10468 14816
rect 11428 14807 11480 14816
rect 11428 14773 11437 14807
rect 11437 14773 11471 14807
rect 11471 14773 11480 14807
rect 11428 14764 11480 14773
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 12808 14764 12860 14816
rect 13636 14807 13688 14816
rect 13636 14773 13645 14807
rect 13645 14773 13679 14807
rect 13679 14773 13688 14807
rect 13636 14764 13688 14773
rect 14096 14807 14148 14816
rect 14096 14773 14105 14807
rect 14105 14773 14139 14807
rect 14139 14773 14148 14807
rect 14096 14764 14148 14773
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 4620 14603 4672 14612
rect 4620 14569 4629 14603
rect 4629 14569 4663 14603
rect 4663 14569 4672 14603
rect 4620 14560 4672 14569
rect 9220 14560 9272 14612
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4528 14356 4580 14408
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 5172 14399 5224 14408
rect 5172 14365 5181 14399
rect 5181 14365 5215 14399
rect 5215 14365 5224 14399
rect 5172 14356 5224 14365
rect 3240 14220 3292 14272
rect 5816 14424 5868 14476
rect 7380 14492 7432 14544
rect 6736 14424 6788 14476
rect 9036 14424 9088 14476
rect 9128 14356 9180 14408
rect 13636 14492 13688 14544
rect 14188 14492 14240 14544
rect 11888 14424 11940 14476
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11244 14356 11296 14408
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 13084 14356 13136 14408
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 10784 14263 10836 14272
rect 10784 14229 10793 14263
rect 10793 14229 10827 14263
rect 10827 14229 10836 14263
rect 10784 14220 10836 14229
rect 11796 14220 11848 14272
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 4528 14059 4580 14068
rect 4528 14025 4537 14059
rect 4537 14025 4571 14059
rect 4571 14025 4580 14059
rect 4528 14016 4580 14025
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 6276 14059 6328 14068
rect 6276 14025 6285 14059
rect 6285 14025 6319 14059
rect 6319 14025 6328 14059
rect 6276 14016 6328 14025
rect 6736 14059 6788 14068
rect 6736 14025 6745 14059
rect 6745 14025 6779 14059
rect 6779 14025 6788 14059
rect 6736 14016 6788 14025
rect 8392 14016 8444 14068
rect 8944 14016 8996 14068
rect 9036 14059 9088 14068
rect 9036 14025 9045 14059
rect 9045 14025 9079 14059
rect 9079 14025 9088 14059
rect 9036 14016 9088 14025
rect 5172 13948 5224 14000
rect 7012 13948 7064 14000
rect 10968 14016 11020 14068
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 11888 14016 11940 14025
rect 11980 14016 12032 14068
rect 12808 14059 12860 14068
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 14188 14059 14240 14068
rect 14188 14025 14197 14059
rect 14197 14025 14231 14059
rect 14231 14025 14240 14059
rect 14188 14016 14240 14025
rect 4436 13812 4488 13864
rect 5632 13880 5684 13932
rect 7656 13880 7708 13932
rect 10508 13948 10560 14000
rect 9496 13880 9548 13932
rect 11244 13880 11296 13932
rect 5264 13744 5316 13796
rect 5540 13744 5592 13796
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 8668 13812 8720 13864
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 10232 13812 10284 13864
rect 10600 13812 10652 13864
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 11796 13855 11848 13864
rect 11796 13821 11805 13855
rect 11805 13821 11839 13855
rect 11839 13821 11848 13855
rect 11796 13812 11848 13821
rect 12900 13812 12952 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 12716 13744 12768 13796
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 6460 13719 6512 13728
rect 6460 13685 6469 13719
rect 6469 13685 6503 13719
rect 6503 13685 6512 13719
rect 6460 13676 6512 13685
rect 7472 13676 7524 13728
rect 8668 13676 8720 13728
rect 10600 13676 10652 13728
rect 11244 13676 11296 13728
rect 12992 13676 13044 13728
rect 13820 13676 13872 13728
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 7472 13472 7524 13524
rect 3240 13404 3292 13456
rect 5724 13404 5776 13456
rect 6920 13404 6972 13456
rect 10968 13472 11020 13524
rect 11244 13472 11296 13524
rect 12900 13472 12952 13524
rect 8852 13404 8904 13456
rect 10048 13404 10100 13456
rect 15108 13404 15160 13456
rect 5172 13336 5224 13388
rect 5264 13336 5316 13388
rect 5540 13379 5592 13388
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 5816 13379 5868 13388
rect 5816 13345 5825 13379
rect 5825 13345 5859 13379
rect 5859 13345 5868 13379
rect 5816 13336 5868 13345
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 9404 13379 9456 13388
rect 9404 13345 9438 13379
rect 9438 13345 9456 13379
rect 9404 13336 9456 13345
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 4988 13200 5040 13252
rect 4804 13132 4856 13184
rect 4896 13132 4948 13184
rect 8944 13200 8996 13252
rect 11888 13336 11940 13388
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13176 13336 13228 13388
rect 13084 13268 13136 13320
rect 6920 13132 6972 13184
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 7564 13132 7616 13141
rect 8852 13175 8904 13184
rect 8852 13141 8861 13175
rect 8861 13141 8895 13175
rect 8895 13141 8904 13175
rect 8852 13132 8904 13141
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 11428 13175 11480 13184
rect 11428 13141 11437 13175
rect 11437 13141 11471 13175
rect 11471 13141 11480 13175
rect 11428 13132 11480 13141
rect 11520 13132 11572 13184
rect 13084 13132 13136 13184
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 5724 12928 5776 12980
rect 6276 12928 6328 12980
rect 7196 12928 7248 12980
rect 9404 12928 9456 12980
rect 13268 12928 13320 12980
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4620 12792 4672 12844
rect 7472 12860 7524 12912
rect 8944 12860 8996 12912
rect 4528 12767 4580 12776
rect 4528 12733 4537 12767
rect 4537 12733 4571 12767
rect 4571 12733 4580 12767
rect 4528 12724 4580 12733
rect 4712 12724 4764 12776
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 5172 12724 5224 12776
rect 6460 12835 6512 12844
rect 6460 12801 6469 12835
rect 6469 12801 6503 12835
rect 6503 12801 6512 12835
rect 6460 12792 6512 12801
rect 6368 12724 6420 12776
rect 8576 12792 8628 12844
rect 9036 12792 9088 12844
rect 9496 12792 9548 12844
rect 10784 12792 10836 12844
rect 11428 12792 11480 12844
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 10416 12724 10468 12776
rect 11888 12724 11940 12776
rect 12348 12767 12400 12776
rect 12348 12733 12357 12767
rect 12357 12733 12391 12767
rect 12391 12733 12400 12767
rect 12348 12724 12400 12733
rect 12716 12724 12768 12776
rect 13084 12724 13136 12776
rect 13268 12724 13320 12776
rect 13912 12767 13964 12776
rect 13912 12733 13921 12767
rect 13921 12733 13955 12767
rect 13955 12733 13964 12767
rect 13912 12724 13964 12733
rect 15108 12724 15160 12776
rect 4436 12699 4488 12708
rect 4436 12665 4445 12699
rect 4445 12665 4479 12699
rect 4479 12665 4488 12699
rect 4436 12656 4488 12665
rect 5356 12656 5408 12708
rect 8300 12656 8352 12708
rect 12164 12656 12216 12708
rect 4712 12631 4764 12640
rect 4712 12597 4721 12631
rect 4721 12597 4755 12631
rect 4755 12597 4764 12631
rect 4712 12588 4764 12597
rect 7012 12588 7064 12640
rect 7564 12588 7616 12640
rect 9036 12588 9088 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 13728 12588 13780 12640
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 8116 12384 8168 12436
rect 8392 12384 8444 12436
rect 8668 12384 8720 12436
rect 11428 12384 11480 12436
rect 11888 12384 11940 12436
rect 7472 12359 7524 12368
rect 7472 12325 7481 12359
rect 7481 12325 7515 12359
rect 7515 12325 7524 12359
rect 7472 12316 7524 12325
rect 3608 12291 3660 12300
rect 3608 12257 3617 12291
rect 3617 12257 3651 12291
rect 3651 12257 3660 12291
rect 3608 12248 3660 12257
rect 4160 12291 4212 12300
rect 4160 12257 4167 12291
rect 4167 12257 4212 12291
rect 4160 12248 4212 12257
rect 4344 12291 4396 12300
rect 4344 12257 4353 12291
rect 4353 12257 4387 12291
rect 4387 12257 4396 12291
rect 4344 12248 4396 12257
rect 4804 12248 4856 12300
rect 4528 12180 4580 12232
rect 5356 12291 5408 12300
rect 5356 12257 5365 12291
rect 5365 12257 5399 12291
rect 5399 12257 5408 12291
rect 5356 12248 5408 12257
rect 5632 12248 5684 12300
rect 5448 12044 5500 12096
rect 6552 12044 6604 12096
rect 7012 12291 7064 12300
rect 7012 12257 7021 12291
rect 7021 12257 7055 12291
rect 7055 12257 7064 12291
rect 7012 12248 7064 12257
rect 7196 12291 7248 12300
rect 7196 12257 7205 12291
rect 7205 12257 7239 12291
rect 7239 12257 7248 12291
rect 7196 12248 7248 12257
rect 7288 12248 7340 12300
rect 7748 12248 7800 12300
rect 12624 12316 12676 12368
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 7564 12180 7616 12232
rect 7932 12223 7984 12232
rect 7932 12189 7941 12223
rect 7941 12189 7975 12223
rect 7975 12189 7984 12223
rect 7932 12180 7984 12189
rect 8116 12180 8168 12232
rect 8392 12291 8444 12300
rect 8392 12257 8401 12291
rect 8401 12257 8435 12291
rect 8435 12257 8444 12291
rect 8392 12248 8444 12257
rect 8484 12248 8536 12300
rect 8300 12112 8352 12164
rect 7748 12044 7800 12096
rect 8208 12044 8260 12096
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 11060 12112 11112 12164
rect 12992 12044 13044 12096
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 4528 11840 4580 11892
rect 5080 11840 5132 11892
rect 7380 11883 7432 11892
rect 7380 11849 7389 11883
rect 7389 11849 7423 11883
rect 7423 11849 7432 11883
rect 7380 11840 7432 11849
rect 8392 11840 8444 11892
rect 8576 11840 8628 11892
rect 4160 11704 4212 11756
rect 4712 11704 4764 11756
rect 4436 11636 4488 11688
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 7656 11568 7708 11620
rect 8484 11568 8536 11620
rect 9036 11636 9088 11688
rect 9588 11679 9640 11688
rect 9588 11645 9597 11679
rect 9597 11645 9631 11679
rect 9631 11645 9640 11679
rect 9588 11636 9640 11645
rect 9772 11679 9824 11688
rect 9772 11645 9781 11679
rect 9781 11645 9815 11679
rect 9815 11645 9824 11679
rect 9772 11636 9824 11645
rect 9864 11679 9916 11688
rect 9864 11645 9873 11679
rect 9873 11645 9907 11679
rect 9907 11645 9916 11679
rect 9864 11636 9916 11645
rect 10048 11636 10100 11688
rect 10140 11679 10192 11688
rect 10140 11645 10149 11679
rect 10149 11645 10183 11679
rect 10183 11645 10192 11679
rect 10140 11636 10192 11645
rect 10692 11636 10744 11688
rect 11152 11772 11204 11824
rect 11428 11704 11480 11756
rect 12348 11840 12400 11892
rect 12716 11883 12768 11892
rect 12716 11849 12725 11883
rect 12725 11849 12759 11883
rect 12759 11849 12768 11883
rect 12716 11840 12768 11849
rect 10508 11568 10560 11620
rect 11060 11568 11112 11620
rect 11152 11568 11204 11620
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 7932 11500 7984 11552
rect 8576 11500 8628 11552
rect 10600 11500 10652 11552
rect 10876 11500 10928 11552
rect 11888 11500 11940 11552
rect 12072 11500 12124 11552
rect 13268 11636 13320 11688
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 12808 11500 12860 11552
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 8208 11296 8260 11348
rect 8760 11296 8812 11348
rect 9588 11339 9640 11348
rect 9588 11305 9597 11339
rect 9597 11305 9631 11339
rect 9631 11305 9640 11339
rect 9588 11296 9640 11305
rect 10048 11296 10100 11348
rect 6276 11228 6328 11280
rect 8576 11228 8628 11280
rect 5724 11160 5776 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 6920 11160 6972 11212
rect 5540 11092 5592 11144
rect 5356 10999 5408 11008
rect 5356 10965 5365 10999
rect 5365 10965 5399 10999
rect 5399 10965 5408 10999
rect 5356 10956 5408 10965
rect 5632 10956 5684 11008
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 11060 11296 11112 11348
rect 11888 11296 11940 11348
rect 13176 11296 13228 11348
rect 11428 11228 11480 11280
rect 8944 11160 8996 11212
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 9312 11092 9364 11144
rect 10232 11160 10284 11212
rect 10968 11203 11020 11212
rect 10968 11169 10977 11203
rect 10977 11169 11011 11203
rect 11011 11169 11020 11203
rect 10968 11160 11020 11169
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 10692 11024 10744 11076
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12624 11160 12676 11212
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 13912 11160 13964 11212
rect 12440 11092 12492 11144
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 12992 11092 13044 11144
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 11888 11024 11940 11076
rect 11980 11024 12032 11076
rect 7288 10956 7340 11008
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 10600 10956 10652 11008
rect 11244 10956 11296 11008
rect 12164 10999 12216 11008
rect 12164 10965 12173 10999
rect 12173 10965 12207 10999
rect 12207 10965 12216 10999
rect 12164 10956 12216 10965
rect 12900 10956 12952 11008
rect 13176 10956 13228 11008
rect 13636 10956 13688 11008
rect 15108 10956 15160 11008
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 5264 10684 5316 10736
rect 6276 10752 6328 10804
rect 7380 10752 7432 10804
rect 9588 10752 9640 10804
rect 11612 10752 11664 10804
rect 12256 10752 12308 10804
rect 12532 10752 12584 10804
rect 12716 10752 12768 10804
rect 12900 10752 12952 10804
rect 5816 10684 5868 10736
rect 9220 10684 9272 10736
rect 7932 10616 7984 10668
rect 8392 10616 8444 10668
rect 10968 10616 11020 10668
rect 5172 10548 5224 10600
rect 4620 10480 4672 10532
rect 5356 10480 5408 10532
rect 5724 10480 5776 10532
rect 4528 10412 4580 10464
rect 4896 10412 4948 10464
rect 5632 10412 5684 10464
rect 8944 10548 8996 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10140 10548 10192 10600
rect 11152 10548 11204 10600
rect 12164 10616 12216 10668
rect 12256 10591 12308 10600
rect 12256 10557 12265 10591
rect 12265 10557 12299 10591
rect 12299 10557 12308 10591
rect 12256 10548 12308 10557
rect 9588 10480 9640 10532
rect 11060 10480 11112 10532
rect 12624 10548 12676 10600
rect 14924 10659 14976 10668
rect 14924 10625 14933 10659
rect 14933 10625 14967 10659
rect 14967 10625 14976 10659
rect 14924 10616 14976 10625
rect 15108 10548 15160 10600
rect 9036 10412 9088 10464
rect 11428 10412 11480 10464
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 12440 10412 12492 10464
rect 14924 10480 14976 10532
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 13084 10412 13136 10464
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 4620 10208 4672 10260
rect 5264 10208 5316 10260
rect 5724 10208 5776 10260
rect 6460 10208 6512 10260
rect 6920 10208 6972 10260
rect 4528 10140 4580 10192
rect 8576 10208 8628 10260
rect 4896 10115 4948 10124
rect 4896 10081 4905 10115
rect 4905 10081 4939 10115
rect 4939 10081 4948 10115
rect 4896 10072 4948 10081
rect 5356 10004 5408 10056
rect 5540 10072 5592 10124
rect 6552 10072 6604 10124
rect 6920 10072 6972 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9404 10208 9456 10260
rect 10140 10208 10192 10260
rect 12992 10208 13044 10260
rect 9128 10072 9180 10124
rect 11244 10183 11296 10192
rect 11244 10149 11253 10183
rect 11253 10149 11287 10183
rect 11287 10149 11296 10183
rect 11244 10140 11296 10149
rect 9496 10115 9548 10124
rect 9496 10081 9530 10115
rect 9530 10081 9548 10115
rect 9496 10072 9548 10081
rect 11152 10072 11204 10124
rect 11796 10183 11848 10192
rect 11796 10149 11805 10183
rect 11805 10149 11839 10183
rect 11839 10149 11848 10183
rect 11796 10140 11848 10149
rect 11888 10140 11940 10192
rect 12532 10140 12584 10192
rect 12900 10140 12952 10192
rect 14924 10140 14976 10192
rect 5632 9936 5684 9988
rect 5816 10004 5868 10056
rect 6644 9936 6696 9988
rect 12164 10072 12216 10124
rect 12808 10072 12860 10124
rect 12992 10115 13044 10124
rect 12992 10081 13001 10115
rect 13001 10081 13035 10115
rect 13035 10081 13044 10115
rect 12992 10072 13044 10081
rect 11980 10004 12032 10056
rect 12716 10004 12768 10056
rect 12256 9936 12308 9988
rect 8392 9868 8444 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 11520 9911 11572 9920
rect 11520 9877 11529 9911
rect 11529 9877 11563 9911
rect 11563 9877 11572 9911
rect 11520 9868 11572 9877
rect 12532 9868 12584 9920
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 5080 9707 5132 9716
rect 5080 9673 5089 9707
rect 5089 9673 5123 9707
rect 5123 9673 5132 9707
rect 5080 9664 5132 9673
rect 6552 9664 6604 9716
rect 11520 9664 11572 9716
rect 5632 9596 5684 9648
rect 5448 9528 5500 9580
rect 8484 9596 8536 9648
rect 5172 9392 5224 9444
rect 5448 9392 5500 9444
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7656 9528 7708 9580
rect 7472 9503 7524 9512
rect 5724 9392 5776 9444
rect 5908 9435 5960 9444
rect 5908 9401 5917 9435
rect 5917 9401 5951 9435
rect 5951 9401 5960 9435
rect 5908 9392 5960 9401
rect 6460 9435 6512 9444
rect 6460 9401 6469 9435
rect 6469 9401 6503 9435
rect 6503 9401 6512 9435
rect 6460 9392 6512 9401
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 8944 9460 8996 9512
rect 15016 9528 15068 9580
rect 7564 9392 7616 9444
rect 10232 9392 10284 9444
rect 11428 9460 11480 9512
rect 12624 9460 12676 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 13084 9460 13136 9512
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 14924 9460 14976 9512
rect 14004 9392 14056 9444
rect 3884 9324 3936 9376
rect 6736 9324 6788 9376
rect 6828 9367 6880 9376
rect 6828 9333 6837 9367
rect 6837 9333 6871 9367
rect 6871 9333 6880 9367
rect 6828 9324 6880 9333
rect 7104 9324 7156 9376
rect 9312 9324 9364 9376
rect 10968 9324 11020 9376
rect 11060 9324 11112 9376
rect 12624 9367 12676 9376
rect 12624 9333 12633 9367
rect 12633 9333 12667 9367
rect 12667 9333 12676 9367
rect 12624 9324 12676 9333
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 5080 9163 5132 9172
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5632 9120 5684 9172
rect 6552 9120 6604 9172
rect 6828 9120 6880 9172
rect 8944 9120 8996 9172
rect 9496 9120 9548 9172
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 3608 9027 3660 9036
rect 3608 8993 3642 9027
rect 3642 8993 3660 9027
rect 3608 8984 3660 8993
rect 5908 9052 5960 9104
rect 6368 9052 6420 9104
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 8760 9052 8812 9104
rect 5540 9027 5592 9036
rect 5540 8993 5549 9027
rect 5549 8993 5583 9027
rect 5583 8993 5592 9027
rect 5540 8984 5592 8993
rect 5724 8984 5776 9036
rect 7012 8984 7064 9036
rect 8852 8984 8904 9036
rect 8944 9027 8996 9036
rect 8944 8993 8953 9027
rect 8953 8993 8987 9027
rect 8987 8993 8996 9027
rect 8944 8984 8996 8993
rect 9036 8984 9088 9036
rect 9220 9027 9272 9036
rect 9220 8993 9229 9027
rect 9229 8993 9263 9027
rect 9263 8993 9272 9027
rect 9220 8984 9272 8993
rect 9404 8984 9456 9036
rect 10324 9052 10376 9104
rect 5448 8916 5500 8968
rect 7288 8916 7340 8968
rect 7472 8916 7524 8968
rect 10692 8984 10744 9036
rect 12808 9052 12860 9104
rect 6920 8891 6972 8900
rect 6920 8857 6929 8891
rect 6929 8857 6963 8891
rect 6963 8857 6972 8891
rect 6920 8848 6972 8857
rect 10600 8916 10652 8968
rect 12440 8984 12492 9036
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 13912 9120 13964 9172
rect 13268 8916 13320 8968
rect 13084 8848 13136 8900
rect 3976 8780 4028 8832
rect 8576 8780 8628 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 3608 8576 3660 8628
rect 5632 8576 5684 8628
rect 6736 8576 6788 8628
rect 3884 8415 3936 8424
rect 3884 8381 3893 8415
rect 3893 8381 3927 8415
rect 3927 8381 3936 8415
rect 3884 8372 3936 8381
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 6460 8415 6512 8424
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 6460 8372 6512 8381
rect 6644 8415 6696 8424
rect 6644 8381 6653 8415
rect 6653 8381 6687 8415
rect 6687 8381 6696 8415
rect 6644 8372 6696 8381
rect 6736 8372 6788 8424
rect 7472 8576 7524 8628
rect 8944 8576 8996 8628
rect 9312 8576 9364 8628
rect 12716 8576 12768 8628
rect 8208 8440 8260 8492
rect 8392 8483 8444 8492
rect 8392 8449 8401 8483
rect 8401 8449 8435 8483
rect 8435 8449 8444 8483
rect 8392 8440 8444 8449
rect 11428 8551 11480 8560
rect 11428 8517 11437 8551
rect 11437 8517 11471 8551
rect 11471 8517 11480 8551
rect 11428 8508 11480 8517
rect 8300 8372 8352 8424
rect 8668 8372 8720 8424
rect 9404 8440 9456 8492
rect 10784 8440 10836 8492
rect 8852 8415 8904 8424
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 7564 8304 7616 8356
rect 9404 8304 9456 8356
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12808 8440 12860 8492
rect 10600 8304 10652 8356
rect 12624 8372 12676 8424
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14924 8372 14976 8424
rect 5816 8236 5868 8288
rect 7104 8236 7156 8288
rect 8944 8236 8996 8288
rect 9036 8279 9088 8288
rect 9036 8245 9045 8279
rect 9045 8245 9079 8279
rect 9079 8245 9088 8279
rect 9036 8236 9088 8245
rect 11152 8236 11204 8288
rect 13084 8304 13136 8356
rect 13176 8236 13228 8288
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 7104 8032 7156 8084
rect 8208 8032 8260 8084
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 9404 8075 9456 8084
rect 9404 8041 9413 8075
rect 9413 8041 9447 8075
rect 9447 8041 9456 8075
rect 9404 8032 9456 8041
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 6460 7896 6512 7948
rect 7104 7896 7156 7948
rect 8300 8007 8352 8016
rect 8300 7973 8309 8007
rect 8309 7973 8343 8007
rect 8343 7973 8352 8007
rect 8300 7964 8352 7973
rect 8760 8007 8812 8016
rect 8760 7973 8795 8007
rect 8795 7973 8812 8007
rect 8760 7964 8812 7973
rect 9036 7964 9088 8016
rect 7564 7760 7616 7812
rect 10416 7939 10468 7948
rect 10416 7905 10425 7939
rect 10425 7905 10459 7939
rect 10459 7905 10468 7939
rect 10416 7896 10468 7905
rect 11428 7896 11480 7948
rect 12900 7828 12952 7880
rect 13268 7828 13320 7880
rect 6276 7692 6328 7744
rect 6828 7692 6880 7744
rect 8208 7692 8260 7744
rect 8484 7735 8536 7744
rect 8484 7701 8493 7735
rect 8493 7701 8527 7735
rect 8527 7701 8536 7735
rect 8484 7692 8536 7701
rect 8944 7735 8996 7744
rect 8944 7701 8953 7735
rect 8953 7701 8987 7735
rect 8987 7701 8996 7735
rect 8944 7692 8996 7701
rect 13728 7692 13780 7744
rect 14740 7735 14792 7744
rect 14740 7701 14749 7735
rect 14749 7701 14783 7735
rect 14783 7701 14792 7735
rect 14740 7692 14792 7701
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 5540 7488 5592 7540
rect 6644 7488 6696 7540
rect 10692 7488 10744 7540
rect 11244 7488 11296 7540
rect 7748 7463 7800 7472
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 10508 7420 10560 7472
rect 12900 7463 12952 7472
rect 12900 7429 12909 7463
rect 12909 7429 12943 7463
rect 12943 7429 12952 7463
rect 12900 7420 12952 7429
rect 5724 7352 5776 7404
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 6368 7327 6420 7336
rect 5632 7284 5684 7293
rect 6368 7293 6377 7327
rect 6377 7293 6411 7327
rect 6411 7293 6420 7327
rect 6368 7284 6420 7293
rect 5816 7216 5868 7268
rect 6460 7216 6512 7268
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 7656 7352 7708 7404
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 7564 7284 7616 7336
rect 8208 7284 8260 7336
rect 11336 7327 11388 7336
rect 11336 7293 11345 7327
rect 11345 7293 11379 7327
rect 11379 7293 11388 7327
rect 11336 7284 11388 7293
rect 12072 7352 12124 7404
rect 5264 7148 5316 7200
rect 6736 7148 6788 7200
rect 7380 7216 7432 7268
rect 10968 7216 11020 7268
rect 13728 7284 13780 7336
rect 11888 7216 11940 7268
rect 11060 7148 11112 7200
rect 11336 7148 11388 7200
rect 12256 7148 12308 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 14004 7191 14056 7200
rect 14004 7157 14013 7191
rect 14013 7157 14047 7191
rect 14047 7157 14056 7191
rect 14004 7148 14056 7157
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 6460 6944 6512 6996
rect 5724 6876 5776 6928
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 5816 6808 5868 6860
rect 6368 6919 6420 6928
rect 6368 6885 6377 6919
rect 6377 6885 6411 6919
rect 6411 6885 6420 6919
rect 6368 6876 6420 6885
rect 8484 6944 8536 6996
rect 4068 6604 4120 6656
rect 5632 6672 5684 6724
rect 5908 6672 5960 6724
rect 5494 6604 5546 6656
rect 6920 6808 6972 6860
rect 7472 6808 7524 6860
rect 7748 6851 7800 6860
rect 7748 6817 7757 6851
rect 7757 6817 7791 6851
rect 7791 6817 7800 6851
rect 7748 6808 7800 6817
rect 8208 6876 8260 6928
rect 8484 6808 8536 6860
rect 12072 6944 12124 6996
rect 11888 6876 11940 6928
rect 6552 6740 6604 6792
rect 7196 6740 7248 6792
rect 7656 6740 7708 6792
rect 8392 6783 8444 6792
rect 8392 6749 8401 6783
rect 8401 6749 8435 6783
rect 8435 6749 8444 6783
rect 8392 6740 8444 6749
rect 6276 6672 6328 6724
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 12440 6808 12492 6860
rect 12900 6851 12952 6860
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 13176 6944 13228 6996
rect 14740 6944 14792 6996
rect 13544 6919 13596 6928
rect 13544 6885 13553 6919
rect 13553 6885 13587 6919
rect 13587 6885 13596 6919
rect 13544 6876 13596 6885
rect 13084 6808 13136 6860
rect 13728 6808 13780 6860
rect 11060 6740 11112 6792
rect 6460 6604 6512 6656
rect 6736 6647 6788 6656
rect 6736 6613 6745 6647
rect 6745 6613 6779 6647
rect 6779 6613 6788 6647
rect 6736 6604 6788 6613
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 12256 6783 12308 6792
rect 12256 6749 12265 6783
rect 12265 6749 12299 6783
rect 12299 6749 12308 6783
rect 12256 6740 12308 6749
rect 12348 6740 12400 6792
rect 12716 6672 12768 6724
rect 12164 6604 12216 6656
rect 12348 6604 12400 6656
rect 12624 6604 12676 6656
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 13084 6604 13136 6613
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 5632 6400 5684 6452
rect 6276 6400 6328 6452
rect 7380 6400 7432 6452
rect 7748 6400 7800 6452
rect 12716 6443 12768 6452
rect 12716 6409 12725 6443
rect 12725 6409 12759 6443
rect 12759 6409 12768 6443
rect 12716 6400 12768 6409
rect 12900 6400 12952 6452
rect 14004 6400 14056 6452
rect 6000 6332 6052 6384
rect 6460 6264 6512 6316
rect 6736 6332 6788 6384
rect 6644 6264 6696 6316
rect 8300 6264 8352 6316
rect 9128 6264 9180 6316
rect 3976 6196 4028 6248
rect 5724 6239 5776 6248
rect 5724 6205 5733 6239
rect 5733 6205 5767 6239
rect 5767 6205 5776 6239
rect 5724 6196 5776 6205
rect 6368 6239 6420 6248
rect 6368 6205 6377 6239
rect 6377 6205 6411 6239
rect 6411 6205 6420 6239
rect 6368 6196 6420 6205
rect 7104 6239 7156 6248
rect 7104 6205 7113 6239
rect 7113 6205 7147 6239
rect 7147 6205 7156 6239
rect 7104 6196 7156 6205
rect 7564 6196 7616 6248
rect 9404 6196 9456 6248
rect 10508 6196 10560 6248
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 4896 6128 4948 6180
rect 6000 6171 6052 6180
rect 6000 6137 6009 6171
rect 6009 6137 6043 6171
rect 6043 6137 6052 6171
rect 6000 6128 6052 6137
rect 6552 6128 6604 6180
rect 10324 6128 10376 6180
rect 14924 6196 14976 6248
rect 5356 6060 5408 6112
rect 11060 6060 11112 6112
rect 12072 6060 12124 6112
rect 12440 6060 12492 6112
rect 12808 6060 12860 6112
rect 13176 6103 13228 6112
rect 13176 6069 13201 6103
rect 13201 6069 13228 6103
rect 13176 6060 13228 6069
rect 13820 6060 13872 6112
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 6000 5720 6052 5772
rect 6276 5720 6328 5772
rect 6644 5788 6696 5840
rect 7380 5788 7432 5840
rect 6736 5720 6788 5772
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8944 5856 8996 5908
rect 8668 5831 8720 5840
rect 8668 5797 8695 5831
rect 8695 5797 8720 5831
rect 8668 5788 8720 5797
rect 8760 5788 8812 5840
rect 10784 5856 10836 5908
rect 11428 5856 11480 5908
rect 11980 5856 12032 5908
rect 10324 5788 10376 5840
rect 5724 5584 5776 5636
rect 6828 5584 6880 5636
rect 10048 5720 10100 5772
rect 12624 5720 12676 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 13176 5763 13228 5772
rect 13176 5729 13185 5763
rect 13185 5729 13219 5763
rect 13219 5729 13228 5763
rect 13176 5720 13228 5729
rect 13268 5720 13320 5772
rect 10140 5627 10192 5636
rect 10140 5593 10149 5627
rect 10149 5593 10183 5627
rect 10183 5593 10192 5627
rect 10140 5584 10192 5593
rect 13084 5652 13136 5704
rect 5172 5516 5224 5568
rect 6920 5516 6972 5568
rect 7012 5516 7064 5568
rect 8300 5516 8352 5568
rect 9312 5516 9364 5568
rect 10232 5516 10284 5568
rect 11060 5516 11112 5568
rect 11796 5516 11848 5568
rect 13084 5516 13136 5568
rect 14924 5559 14976 5568
rect 14924 5525 14933 5559
rect 14933 5525 14967 5559
rect 14967 5525 14976 5559
rect 14924 5516 14976 5525
rect 15660 5516 15712 5568
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 4896 5355 4948 5364
rect 4896 5321 4905 5355
rect 4905 5321 4939 5355
rect 4939 5321 4948 5355
rect 4896 5312 4948 5321
rect 10324 5312 10376 5364
rect 11244 5312 11296 5364
rect 5816 5244 5868 5296
rect 7104 5244 7156 5296
rect 8208 5244 8260 5296
rect 10140 5244 10192 5296
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 5356 5151 5408 5160
rect 5356 5117 5365 5151
rect 5365 5117 5399 5151
rect 5399 5117 5408 5151
rect 5356 5108 5408 5117
rect 5724 5108 5776 5160
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 6276 5219 6328 5228
rect 6276 5185 6285 5219
rect 6285 5185 6319 5219
rect 6319 5185 6328 5219
rect 6276 5176 6328 5185
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7748 5176 7800 5228
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 10048 5176 10100 5228
rect 6368 5108 6420 5160
rect 6828 5108 6880 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7104 5108 7156 5160
rect 8300 5108 8352 5160
rect 6000 5040 6052 5092
rect 9772 5040 9824 5092
rect 10232 5040 10284 5092
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 11796 5219 11848 5228
rect 11796 5185 11805 5219
rect 11805 5185 11839 5219
rect 11839 5185 11848 5219
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 12992 5312 13044 5364
rect 12900 5244 12952 5296
rect 11796 5176 11848 5185
rect 11428 5151 11480 5160
rect 11428 5117 11437 5151
rect 11437 5117 11471 5151
rect 11471 5117 11480 5151
rect 11428 5108 11480 5117
rect 13176 5176 13228 5228
rect 14648 5176 14700 5228
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 7472 5015 7524 5024
rect 7472 4981 7481 5015
rect 7481 4981 7515 5015
rect 7515 4981 7524 5015
rect 7472 4972 7524 4981
rect 10324 5015 10376 5024
rect 10324 4981 10333 5015
rect 10333 4981 10367 5015
rect 10367 4981 10376 5015
rect 10324 4972 10376 4981
rect 10508 4972 10560 5024
rect 11888 5040 11940 5092
rect 12440 5108 12492 5160
rect 13728 5040 13780 5092
rect 12072 4972 12124 5024
rect 12164 5015 12216 5024
rect 12164 4981 12173 5015
rect 12173 4981 12207 5015
rect 12207 4981 12216 5015
rect 12164 4972 12216 4981
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 5724 4768 5776 4820
rect 6000 4768 6052 4820
rect 6276 4768 6328 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 8668 4811 8720 4820
rect 8668 4777 8677 4811
rect 8677 4777 8711 4811
rect 8711 4777 8720 4811
rect 8668 4768 8720 4777
rect 9312 4768 9364 4820
rect 9680 4768 9732 4820
rect 10416 4768 10468 4820
rect 7472 4700 7524 4752
rect 11888 4768 11940 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 3976 4632 4028 4684
rect 4344 4675 4396 4684
rect 4344 4641 4378 4675
rect 4378 4641 4396 4675
rect 4344 4632 4396 4641
rect 6000 4675 6052 4684
rect 6000 4641 6009 4675
rect 6009 4641 6043 4675
rect 6043 4641 6052 4675
rect 6000 4632 6052 4641
rect 6460 4632 6512 4684
rect 7104 4632 7156 4684
rect 8392 4632 8444 4684
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9128 4632 9180 4684
rect 10232 4632 10284 4684
rect 10508 4632 10560 4684
rect 11060 4632 11112 4684
rect 11244 4632 11296 4684
rect 12164 4700 12216 4752
rect 13084 4700 13136 4752
rect 8208 4564 8260 4616
rect 9680 4607 9732 4616
rect 9680 4573 9689 4607
rect 9689 4573 9723 4607
rect 9723 4573 9732 4607
rect 9680 4564 9732 4573
rect 9772 4607 9824 4616
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 10140 4564 10192 4616
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 12072 4496 12124 4548
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 10232 4471 10284 4480
rect 10232 4437 10241 4471
rect 10241 4437 10275 4471
rect 10275 4437 10284 4471
rect 10232 4428 10284 4437
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 4344 4224 4396 4276
rect 5816 4224 5868 4276
rect 6276 4224 6328 4276
rect 10232 4267 10284 4276
rect 10232 4233 10241 4267
rect 10241 4233 10275 4267
rect 10275 4233 10284 4267
rect 10232 4224 10284 4233
rect 8760 4020 8812 4072
rect 5724 3952 5776 4004
rect 6460 3952 6512 4004
rect 10324 3952 10376 4004
rect 5632 3884 5684 3936
rect 6368 3884 6420 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 10508 3680 10560 3732
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 10048 3544 10100 3596
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 10048 3179 10100 3188
rect 10048 3145 10057 3179
rect 10057 3145 10091 3179
rect 10091 3145 10100 3179
rect 10048 3136 10100 3145
rect 10416 2932 10468 2984
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
<< metal2 >>
rect 846 15722 902 16000
rect 846 15694 980 15722
rect 846 15600 902 15694
rect 952 15026 980 15694
rect 2134 15600 2190 16000
rect 3422 15722 3478 16000
rect 4710 15722 4766 16000
rect 3422 15694 3556 15722
rect 3422 15600 3478 15694
rect 940 15020 992 15026
rect 940 14962 992 14968
rect 2148 14958 2176 15600
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 3528 14958 3556 15694
rect 4710 15694 4844 15722
rect 4710 15600 4766 15694
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 2136 14952 2188 14958
rect 2136 14894 2188 14900
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 14278 3280 14350
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 3252 13462 3280 14214
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 3620 12306 3648 14758
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 4448 13870 4476 14962
rect 4816 14958 4844 15694
rect 5998 15600 6054 16000
rect 7286 15600 7342 16000
rect 8574 15722 8630 16000
rect 8574 15694 8708 15722
rect 8574 15600 8630 15694
rect 6012 15450 6040 15600
rect 5828 15422 6040 15450
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4632 14618 4660 14894
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4540 14074 4568 14350
rect 4724 14074 4752 14758
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4160 12776 4212 12782
rect 3988 12724 4160 12730
rect 3988 12718 4212 12724
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 3988 12702 4200 12718
rect 4436 12708 4488 12714
rect 3988 12434 4016 12702
rect 4436 12650 4488 12656
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 3988 12406 4200 12434
rect 4172 12306 4200 12406
rect 4448 12322 4476 12650
rect 4356 12306 4476 12322
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4344 12300 4476 12306
rect 4396 12294 4476 12300
rect 4344 12242 4396 12248
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 4172 11762 4200 12242
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4448 11694 4476 12294
rect 4540 12238 4568 12718
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11898 4568 12174
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4632 11694 4660 12786
rect 4724 12782 4752 14010
rect 5000 13258 5028 14758
rect 5092 14414 5120 15030
rect 5828 14958 5856 15422
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 7300 14958 7328 15600
rect 8680 14958 8708 15694
rect 9862 15600 9918 16000
rect 11150 15600 11206 16000
rect 12438 15600 12494 16000
rect 13726 15600 13782 16000
rect 15014 15600 15070 16000
rect 9876 15450 9904 15600
rect 9876 15422 10088 15450
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 10060 14958 10088 15422
rect 11164 14958 11192 15600
rect 12452 14958 12480 15600
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 13740 14958 13768 15600
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 11152 14952 11204 14958
rect 11152 14894 11204 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 4988 13252 5040 13258
rect 4988 13194 5040 13200
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4816 12782 4844 13126
rect 4908 12986 4936 13126
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4724 11762 4752 12582
rect 4816 12306 4844 12718
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 5092 11898 5120 14350
rect 5184 14006 5212 14350
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5184 13394 5212 13942
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 5540 13796 5592 13802
rect 5644 13784 5672 13874
rect 5592 13756 5672 13784
rect 5540 13738 5592 13744
rect 5276 13394 5304 13738
rect 5552 13394 5580 13738
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5184 12782 5212 13330
rect 5736 12986 5764 13398
rect 5828 13394 5856 14418
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 6276 14068 6328 14074
rect 6276 14010 6328 14016
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12306 5396 12650
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5080 11892 5132 11898
rect 5080 11834 5132 11840
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4436 11688 4488 11694
rect 4436 11630 4488 11636
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 4540 10470 4568 11630
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 4540 10198 4568 10406
rect 4632 10266 4660 10474
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4908 10130 4936 10406
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 3620 8634 3648 8978
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3896 8430 3924 9318
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 5092 9178 5120 9658
rect 5184 9450 5212 10542
rect 5276 10266 5304 10678
rect 5368 10538 5396 10950
rect 5356 10532 5408 10538
rect 5356 10474 5408 10480
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5368 10062 5396 10474
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5460 9586 5488 12038
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5552 10248 5580 11086
rect 5644 11014 5672 12242
rect 5828 11218 5856 13330
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 6288 12986 6316 14010
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6380 12782 6408 14758
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6748 14074 6776 14418
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6932 13870 6960 14758
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7024 13870 7052 13942
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 12850 6500 13670
rect 6932 13462 6960 13806
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6932 12782 6960 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10470 5672 10950
rect 5736 10538 5764 11154
rect 5828 10742 5856 11154
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 6288 10810 6316 11222
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5736 10266 5764 10474
rect 5724 10260 5776 10266
rect 5552 10220 5672 10248
rect 5644 10146 5672 10220
rect 5724 10202 5776 10208
rect 5540 10124 5592 10130
rect 5644 10118 5764 10146
rect 5540 10066 5592 10072
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5460 8974 5488 9386
rect 5552 9042 5580 10066
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5644 9654 5672 9930
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5644 9518 5672 9590
rect 5736 9568 5764 10118
rect 5828 10062 5856 10678
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 5736 9540 5856 9568
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 8430 4016 8774
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 3988 6644 4016 8366
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 5552 7546 5580 8978
rect 5644 8634 5672 9114
rect 5736 9042 5764 9386
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5828 8378 5856 9540
rect 6472 9450 6500 10202
rect 6564 10130 6592 12038
rect 6932 11218 6960 12718
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12306 7052 12582
rect 7208 12306 7236 12922
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7300 11014 7328 12242
rect 7392 11898 7420 14486
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7484 13530 7512 13670
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 13190 7604 14214
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7668 13394 7696 13874
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7484 12374 7512 12854
rect 7576 12646 7604 13126
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 7564 12640 7616 12646
rect 7564 12582 7616 12588
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7576 12238 7604 12582
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 7654 12336 7710 12345
rect 7654 12271 7710 12280
rect 7748 12300 7800 12306
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7668 11626 7696 12271
rect 7748 12242 7800 12248
rect 7760 12102 7788 12242
rect 8128 12238 8156 12378
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6920 10260 6972 10266
rect 7300 10248 7328 10950
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 6972 10220 7328 10248
rect 6920 10202 6972 10208
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6564 9722 6592 10066
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 6460 9444 6512 9450
rect 6460 9386 6512 9392
rect 5920 9110 5948 9386
rect 6472 9330 6500 9386
rect 6380 9302 6500 9330
rect 6380 9110 6408 9302
rect 6564 9178 6592 9658
rect 6552 9172 6604 9178
rect 6472 9132 6552 9160
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 6472 8430 6500 9132
rect 6552 9114 6604 9120
rect 6656 8514 6684 9930
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6748 8634 6776 9318
rect 6840 9178 6868 9318
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 8906 6960 10066
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 7024 9042 7052 9454
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6656 8486 6776 8514
rect 6748 8430 6776 8486
rect 5736 8350 5856 8378
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6644 8424 6696 8430
rect 6644 8366 6696 8372
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5736 7410 5764 8350
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 5276 6866 5304 7142
rect 5644 7018 5672 7278
rect 5506 6990 5672 7018
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5506 6662 5534 6990
rect 5736 6934 5764 7346
rect 5828 7274 5856 8230
rect 6472 7954 6500 8366
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5722 6760 5778 6769
rect 5632 6724 5684 6730
rect 5722 6695 5778 6704
rect 5632 6666 5684 6672
rect 4068 6656 4120 6662
rect 3988 6616 4068 6644
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 3988 6254 4016 6616
rect 4068 6598 4120 6604
rect 5494 6656 5546 6662
rect 5494 6598 5546 6604
rect 5644 6458 5672 6666
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 6254 5764 6695
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 3988 4690 4016 6190
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 4908 5370 4936 6122
rect 5356 6112 5408 6118
rect 5828 6100 5856 6802
rect 5906 6760 5962 6769
rect 6288 6730 6316 7686
rect 6656 7546 6684 8366
rect 7116 8294 7144 9318
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7300 8974 7328 9046
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 7116 8090 7144 8230
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6840 7342 6868 7686
rect 7116 7410 7144 7890
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6380 6934 6408 7278
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6472 7002 6500 7210
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6472 6746 6500 6938
rect 5906 6695 5908 6704
rect 5960 6695 5962 6704
rect 6276 6724 6328 6730
rect 5908 6666 5960 6672
rect 6276 6666 6328 6672
rect 6380 6718 6500 6746
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 6288 6458 6316 6666
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 6012 6186 6040 6326
rect 6380 6254 6408 6718
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6322 6500 6598
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5356 6054 5408 6060
rect 5736 6072 5856 6100
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5184 5166 5212 5510
rect 5368 5166 5396 6054
rect 5736 5642 5764 6072
rect 6012 5778 6040 6122
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5736 5166 5764 5578
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5828 5166 5856 5238
rect 6288 5234 6316 5714
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6380 5166 6408 6190
rect 6564 6186 6592 6734
rect 6748 6662 6776 7142
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6390 6776 6598
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6552 6180 6604 6186
rect 6552 6122 6604 6128
rect 6656 5846 6684 6258
rect 6644 5840 6696 5846
rect 6644 5782 6696 5788
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 4356 4282 4384 4626
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 5644 3942 5672 4966
rect 6012 4826 6040 5034
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 6276 4820 6328 4826
rect 6276 4762 6328 4768
rect 5736 4010 5764 4762
rect 6012 4690 6040 4762
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5828 4282 5856 4422
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 6288 4282 6316 4762
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 6380 3942 6408 5102
rect 6748 4826 6776 5714
rect 6932 5658 6960 6802
rect 7208 6798 7236 7346
rect 7392 7274 7420 10746
rect 7668 9586 7696 11562
rect 7944 11558 7972 12174
rect 8220 12102 8248 12242
rect 8312 12170 8340 12650
rect 8404 12442 8432 14010
rect 8864 13870 8892 14758
rect 8956 14074 8984 14758
rect 9232 14618 9260 14894
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9048 14074 9076 14418
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8680 13734 8708 13806
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13394 8708 13670
rect 8852 13456 8904 13462
rect 8852 13398 8904 13404
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8864 13190 8892 13398
rect 9140 13326 9168 14350
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8956 12918 8984 13194
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 9048 12850 9076 13126
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 8220 11354 8248 12038
rect 8404 11898 8432 12242
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8496 11626 8524 12242
rect 8588 11898 8616 12786
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8588 11286 8616 11494
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7944 10674 7972 10950
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 8404 9926 8432 10610
rect 8588 10266 8616 11222
rect 8680 11218 8708 12378
rect 9048 11694 9076 12582
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8772 11354 8800 11630
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 10606 8984 11154
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8576 10260 8628 10266
rect 8496 10220 8576 10248
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 8974 7512 9454
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7392 6458 7420 7210
rect 7484 6866 7512 8570
rect 7576 8362 7604 9386
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 7818 7604 8298
rect 7668 8022 7696 9522
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 8404 8498 8432 9862
rect 8496 9654 8524 10220
rect 8576 10202 8628 10208
rect 8956 10130 8984 10542
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8588 8838 8616 9862
rect 8956 9518 8984 10066
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8956 9178 8984 9454
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8942 9072 8998 9081
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 8220 8090 8248 8434
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7564 7812 7616 7818
rect 7564 7754 7616 7760
rect 7576 7342 7604 7754
rect 7668 7410 7696 7958
rect 8220 7750 8248 8026
rect 8312 8022 8340 8366
rect 8300 8016 8352 8022
rect 8300 7958 8352 7964
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 6840 5642 6960 5658
rect 6828 5636 6960 5642
rect 6880 5630 6960 5636
rect 6828 5578 6880 5584
rect 6840 5166 6868 5578
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6932 5166 6960 5510
rect 7024 5234 7052 5510
rect 7116 5302 7144 6190
rect 7392 5846 7420 6394
rect 7576 6254 7604 7278
rect 7760 7188 7788 7414
rect 8220 7342 8248 7686
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 7668 7160 7788 7188
rect 7668 6798 7696 7160
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 8220 6934 8248 7278
rect 8208 6928 8260 6934
rect 8404 6882 8432 8434
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 8090 8708 8366
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8772 8022 8800 9046
rect 8852 9036 8904 9042
rect 9048 9042 9076 10406
rect 9140 10130 9168 13262
rect 9416 12986 9444 13330
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 12850 9536 13874
rect 10232 13864 10284 13870
rect 10284 13812 10364 13818
rect 10232 13806 10364 13812
rect 10244 13790 10364 13806
rect 10048 13456 10100 13462
rect 10048 13398 10100 13404
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 10060 11694 10088 13398
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10140 11688 10192 11694
rect 10140 11630 10192 11636
rect 9600 11354 9628 11630
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9784 11218 9812 11630
rect 9876 11218 9904 11630
rect 10060 11354 10088 11630
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9232 9042 9260 10678
rect 9324 9382 9352 11086
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9416 10266 9444 10542
rect 9600 10538 9628 10746
rect 10152 10606 10180 11630
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 10152 10266 10180 10542
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8942 9007 8944 9016
rect 8852 8978 8904 8984
rect 8996 9007 8998 9016
rect 9036 9036 9088 9042
rect 8944 8978 8996 8984
rect 9036 8978 9088 8984
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 8864 8430 8892 8978
rect 8956 8634 8984 8978
rect 9324 8634 9352 9318
rect 9416 9042 9444 10202
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9178 9536 10066
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 10244 9450 10272 11154
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 10336 9110 10364 13790
rect 10428 12782 10456 14758
rect 11440 14414 11468 14758
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 11244 14408 11296 14414
rect 11428 14408 11480 14414
rect 11244 14350 11296 14356
rect 11348 14368 11428 14396
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10508 14000 10560 14006
rect 10508 13942 10560 13948
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9416 8498 9444 8978
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 9036 8288 9088 8294
rect 9036 8230 9088 8236
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7002 8524 7686
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8208 6870 8260 6876
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 8312 6854 8432 6882
rect 8496 6866 8524 6938
rect 8484 6860 8536 6866
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7760 6458 7788 6802
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 8312 6322 8340 6854
rect 8484 6802 8536 6808
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7104 5296 7156 5302
rect 7104 5238 7156 5244
rect 7760 5234 7788 5714
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7104 5160 7156 5166
rect 8220 5137 8248 5238
rect 8312 5166 8340 5510
rect 8404 5234 8432 6734
rect 8772 5846 8800 7958
rect 8956 7750 8984 8230
rect 9048 8022 9076 8230
rect 9416 8090 9444 8298
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 10428 7954 10456 12718
rect 10520 11626 10548 13942
rect 10796 13870 10824 14214
rect 10980 14074 11008 14350
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11256 13938 11284 14350
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10612 13734 10640 13806
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 13530 11284 13670
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10508 11620 10560 11626
rect 10508 11562 10560 11568
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11014 10640 11494
rect 10704 11082 10732 11630
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10169 10640 10950
rect 10598 10160 10654 10169
rect 10598 10095 10654 10104
rect 10612 8974 10640 10095
rect 10704 9178 10732 11018
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10704 9042 10732 9114
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 8944 7744 8996 7750
rect 8944 7686 8996 7692
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 10520 7478 10548 8366
rect 10612 8362 10640 8910
rect 10600 8356 10652 8362
rect 10600 8298 10652 8304
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 5160 8352 5166
rect 7104 5102 7156 5108
rect 8206 5128 8262 5137
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 7116 4690 7144 5102
rect 8300 5102 8352 5108
rect 8206 5063 8262 5072
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4758 7512 4966
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 6472 4010 6500 4626
rect 8220 4622 8248 5063
rect 8404 4690 8432 5170
rect 8680 4826 8708 5782
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8772 4078 8800 5782
rect 8956 4690 8984 5850
rect 9140 5681 9168 6258
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9126 5672 9182 5681
rect 9126 5607 9182 5616
rect 9140 4690 9168 5607
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 4826 9352 5510
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 9416 3602 9444 6190
rect 10336 6186 10364 6598
rect 10520 6254 10548 7414
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 10060 5234 10088 5714
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 10152 5302 10180 5578
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9692 4622 9720 4762
rect 9784 4622 9812 5034
rect 10152 4622 10180 5238
rect 10244 5098 10272 5510
rect 10336 5370 10364 5782
rect 10612 5534 10640 8298
rect 10704 7546 10732 8978
rect 10796 8498 10824 12786
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11098 10916 11494
rect 10980 11218 11008 13466
rect 11060 12164 11112 12170
rect 11060 12106 11112 12112
rect 11072 11626 11100 12106
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11164 11626 11192 11766
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11072 11354 11100 11562
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11218 11192 11562
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11256 11098 11284 13466
rect 10888 11070 11008 11098
rect 10980 10674 11008 11070
rect 11164 11070 11284 11098
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 9382 11008 10610
rect 11164 10606 11192 11070
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10010 11100 10474
rect 11164 10130 11192 10542
rect 11256 10198 11284 10950
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11072 9982 11192 10010
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10796 5914 10824 8434
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10980 5681 11008 7210
rect 11072 7206 11100 9318
rect 11164 8294 11192 9982
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6118 11100 6734
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 10520 5506 10640 5534
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10336 5114 10364 5306
rect 10520 5166 10548 5506
rect 10980 5234 11008 5607
rect 11072 5574 11100 6054
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10508 5160 10560 5166
rect 10506 5128 10508 5137
rect 10560 5128 10562 5137
rect 10232 5092 10284 5098
rect 10336 5086 10456 5114
rect 10232 5034 10284 5040
rect 10244 4690 10272 5034
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 10244 4282 10272 4422
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10336 4010 10364 4966
rect 10428 4826 10456 5086
rect 10506 5063 10562 5072
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10520 4690 10548 4966
rect 11072 4690 11100 5510
rect 11256 5370 11284 7482
rect 11348 7342 11376 14368
rect 11428 14350 11480 14356
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13870 11836 14214
rect 11900 14074 11928 14418
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11796 13864 11848 13870
rect 11848 13824 11928 13852
rect 11796 13806 11848 13812
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 11900 13394 11928 13824
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11440 12850 11468 13126
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11532 12628 11560 13126
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11440 12600 11560 12628
rect 11440 12442 11468 12600
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 11900 12442 11928 12718
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11794 12336 11850 12345
rect 11794 12271 11796 12280
rect 11848 12271 11850 12280
rect 11796 12242 11848 12248
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11286 11468 11698
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 11900 11354 11928 11494
rect 11888 11348 11940 11354
rect 11888 11290 11940 11296
rect 11428 11280 11480 11286
rect 11992 11234 12020 14010
rect 12728 13802 12756 14758
rect 12820 14074 12848 14758
rect 13188 14618 13216 14894
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 14096 14816 14148 14822
rect 14096 14758 14148 14764
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13648 14550 13676 14758
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12912 13530 12940 13806
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 13004 13394 13032 13670
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 13096 13326 13124 14350
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 14108 13870 14136 14758
rect 14188 14544 14240 14550
rect 14188 14486 14240 14492
rect 14200 14074 14228 14486
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13084 13320 13136 13326
rect 13004 13268 13084 13274
rect 13004 13262 13136 13268
rect 13004 13246 13124 13262
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12176 11694 12204 12650
rect 12360 11898 12388 12718
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12374 12664 12582
rect 12624 12368 12676 12374
rect 12624 12310 12676 12316
rect 12728 11898 12756 12718
rect 13004 12102 13032 13246
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12782 13124 13126
rect 13084 12776 13136 12782
rect 13084 12718 13136 12724
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12164 11688 12216 11694
rect 12216 11648 12296 11676
rect 12164 11630 12216 11636
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11428 11222 11480 11228
rect 11900 11206 12020 11234
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10810 11652 11086
rect 11900 11082 11928 11206
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11440 9518 11468 10406
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 11900 10198 11928 10406
rect 11796 10192 11848 10198
rect 11794 10160 11796 10169
rect 11888 10192 11940 10198
rect 11848 10160 11850 10169
rect 11888 10134 11940 10140
rect 11794 10095 11850 10104
rect 11992 10062 12020 11018
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11532 9722 11560 9862
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11440 7954 11468 8502
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 11900 7274 11928 8774
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6866 11376 7142
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 11900 6934 11928 7210
rect 11888 6928 11940 6934
rect 11888 6870 11940 6876
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 11992 5914 12020 9007
rect 12084 7410 12112 11494
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10674 12204 10950
rect 12268 10810 12296 11648
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12440 11144 12492 11150
rect 12346 11112 12402 11121
rect 12440 11086 12492 11092
rect 12346 11047 12402 11056
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12084 7002 12112 7346
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6118 12112 6734
rect 12176 6662 12204 10066
rect 12268 9994 12296 10542
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12360 8498 12388 11047
rect 12452 10470 12480 11086
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12438 10296 12494 10305
rect 12438 10231 12494 10240
rect 12452 9081 12480 10231
rect 12544 10198 12572 10746
rect 12636 10690 12664 11154
rect 12728 10810 12756 11834
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 11218 12848 11494
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 13004 11150 13032 12038
rect 13188 11354 13216 13330
rect 13280 12986 13308 13806
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13355 13084 13663 13093
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13268 12776 13320 12782
rect 13266 12744 13268 12753
rect 13320 12744 13322 12753
rect 13266 12679 13322 12688
rect 13280 11694 13308 12679
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 13740 11694 13768 12582
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13636 11144 13688 11150
rect 13832 11121 13860 13670
rect 13912 12776 13964 12782
rect 13912 12718 13964 12724
rect 13924 11218 13952 12718
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13636 11086 13688 11092
rect 13818 11112 13874 11121
rect 12912 11014 12940 11086
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12636 10662 12848 10690
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9364 12572 9862
rect 12636 9518 12664 10542
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10062 12756 10406
rect 12820 10305 12848 10662
rect 12806 10296 12862 10305
rect 12806 10231 12862 10240
rect 12912 10198 12940 10746
rect 13004 10266 13032 11086
rect 13648 11014 13676 11086
rect 13818 11047 13874 11056
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13004 10130 13032 10202
rect 12808 10124 12860 10130
rect 12808 10066 12860 10072
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12820 9518 12848 10066
rect 13096 9518 13124 10406
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 12624 9376 12676 9382
rect 12544 9336 12624 9364
rect 12624 9318 12676 9324
rect 12438 9072 12494 9081
rect 12438 9007 12440 9016
rect 12492 9007 12494 9016
rect 12440 8978 12492 8984
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12636 8430 12664 9318
rect 12820 9110 12848 9454
rect 13188 9364 13216 10950
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 14922 10704 14978 10713
rect 14922 10639 14924 10648
rect 14976 10639 14978 10648
rect 14924 10610 14976 10616
rect 14936 10538 14964 10610
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 14936 10198 14964 10474
rect 14924 10192 14976 10198
rect 14924 10134 14976 10140
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 15028 9586 15056 15600
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 15106 14512 15162 14521
rect 15106 14447 15162 14456
rect 15120 13462 15148 14447
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 15120 12782 15148 13398
rect 15108 12776 15160 12782
rect 15108 12718 15160 12724
rect 15474 12744 15530 12753
rect 15530 12702 15700 12730
rect 15474 12679 15530 12688
rect 15672 12617 15700 12702
rect 15658 12608 15714 12617
rect 15206 12540 15514 12549
rect 15658 12543 15714 12552
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 15206 11452 15514 11461
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10606 15148 10950
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 13096 9336 13216 9364
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12716 9036 12768 9042
rect 12716 8978 12768 8984
rect 12728 8634 12756 8978
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12820 8498 12848 9046
rect 13096 8906 13124 9336
rect 13924 9178 13952 9454
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13912 9172 13964 9178
rect 13912 9114 13964 9120
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 13096 8362 13124 8842
rect 13084 8356 13136 8362
rect 13084 8298 13136 8304
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7478 12940 7822
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6798 12296 7142
rect 13096 6866 13124 8298
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7002 13216 8230
rect 13280 7886 13308 8910
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 14016 8430 14044 9386
rect 14936 8838 14964 9454
rect 14924 8832 14976 8838
rect 15120 8809 15148 10542
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 14924 8774 14976 8780
rect 15106 8800 15162 8809
rect 14936 8430 14964 8774
rect 15106 8735 15162 8744
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12360 6662 12388 6734
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12452 6254 12480 6802
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12072 6112 12124 6118
rect 12072 6054 12124 6060
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11256 4690 11284 5306
rect 11440 5166 11468 5850
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5234 11836 5510
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 12452 5166 12480 6054
rect 12636 5778 12664 6598
rect 12728 6458 12756 6666
rect 12912 6458 12940 6802
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12820 5370 12848 6054
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12912 5302 12940 6394
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5370 13032 5714
rect 13096 5710 13124 6598
rect 13188 6118 13216 6938
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 13280 5778 13308 7822
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 13740 7342 13768 7686
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 14016 7206 14044 8366
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 13556 6934 13584 7142
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 13176 5772 13228 5778
rect 13176 5714 13228 5720
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12900 5296 12952 5302
rect 12900 5238 12952 5244
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 11900 4826 11928 5034
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 11060 4684 11112 4690
rect 11060 4626 11112 4632
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 10060 3194 10088 3538
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10428 2990 10456 3878
rect 10520 3738 10548 4626
rect 12084 4554 12112 4966
rect 12176 4758 12204 4966
rect 13096 4758 13124 5510
rect 13188 5234 13216 5714
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 13084 4752 13136 4758
rect 13084 4694 13136 4700
rect 13280 4690 13308 5714
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 13740 5098 13768 6802
rect 14016 6458 14044 7142
rect 14752 7002 14780 7686
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14936 6905 14964 8366
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 14922 6896 14978 6905
rect 14922 6831 14978 6840
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 13832 1193 13860 6054
rect 14936 5574 14964 6190
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 15660 5568 15712 5574
rect 15660 5510 15712 5516
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 4826 14688 5170
rect 15672 5001 15700 5510
rect 15658 4992 15714 5001
rect 15206 4924 15514 4933
rect 15658 4927 15714 4936
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14660 4154 14688 4762
rect 14660 4126 14872 4154
rect 14844 3097 14872 4126
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 13818 1184 13874 1193
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 13355 1116 13663 1125
rect 13818 1119 13874 1128
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 7654 12280 7710 12336
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 5722 6704 5778 6760
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 5906 6724 5962 6760
rect 5906 6704 5908 6724
rect 5908 6704 5960 6724
rect 5960 6704 5962 6724
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 8942 9036 8998 9072
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 8942 9016 8944 9036
rect 8944 9016 8996 9036
rect 8996 9016 8998 9036
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 10598 10104 10654 10160
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 8206 5072 8262 5128
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 9126 5616 9182 5672
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 10966 5616 11022 5672
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 10506 5108 10508 5128
rect 10508 5108 10560 5128
rect 10560 5108 10562 5128
rect 10506 5072 10562 5108
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 11794 12300 11850 12336
rect 11794 12280 11796 12300
rect 11796 12280 11848 12300
rect 11848 12280 11850 12300
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 11794 10140 11796 10160
rect 11796 10140 11848 10160
rect 11848 10140 11850 10160
rect 11794 10104 11850 10140
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 11978 9016 12034 9072
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 12346 11056 12402 11112
rect 12438 10240 12494 10296
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 13266 12724 13268 12744
rect 13268 12724 13320 12744
rect 13320 12724 13322 12744
rect 13266 12688 13322 12724
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 12806 10240 12862 10296
rect 13818 11056 13874 11112
rect 12438 9036 12494 9072
rect 12438 9016 12440 9036
rect 12440 9016 12492 9036
rect 12492 9016 12494 9036
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 14922 10668 14978 10704
rect 14922 10648 14924 10668
rect 14924 10648 14976 10668
rect 14976 10648 14978 10668
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 15106 14456 15162 14512
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 15474 12688 15530 12744
rect 15658 12552 15714 12608
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 15106 8744 15162 8800
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 14922 6840 14978 6896
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 15658 4936 15714 4992
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 14830 3032 14886 3088
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 13818 1128 13874 1184
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 15101 14514 15167 14517
rect 15600 14514 16000 14544
rect 15101 14512 16000 14514
rect 15101 14456 15106 14512
rect 15162 14456 16000 14512
rect 15101 14454 16000 14456
rect 15101 14451 15167 14454
rect 15600 14424 16000 14454
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 13351 13023 13667 13024
rect 13261 12746 13327 12749
rect 15469 12746 15535 12749
rect 13261 12744 15535 12746
rect 13261 12688 13266 12744
rect 13322 12688 15474 12744
rect 15530 12688 15535 12744
rect 13261 12686 15535 12688
rect 13261 12683 13327 12686
rect 15469 12683 15535 12686
rect 15600 12608 16000 12640
rect 15600 12552 15658 12608
rect 15714 12552 16000 12608
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15600 12520 16000 12552
rect 15202 12479 15518 12480
rect 7649 12338 7715 12341
rect 11789 12338 11855 12341
rect 7649 12336 11855 12338
rect 7649 12280 7654 12336
rect 7710 12280 11794 12336
rect 11850 12280 11855 12336
rect 7649 12278 11855 12280
rect 7649 12275 7715 12278
rect 11789 12275 11855 12278
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15202 11391 15518 11392
rect 12341 11114 12407 11117
rect 13813 11114 13879 11117
rect 12341 11112 13879 11114
rect 12341 11056 12346 11112
rect 12402 11056 13818 11112
rect 13874 11056 13879 11112
rect 12341 11054 13879 11056
rect 12341 11051 12407 11054
rect 13813 11051 13879 11054
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 14917 10706 14983 10709
rect 15600 10706 16000 10736
rect 14917 10704 16000 10706
rect 14917 10648 14922 10704
rect 14978 10648 16000 10704
rect 14917 10646 16000 10648
rect 14917 10643 14983 10646
rect 15600 10616 16000 10646
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 12433 10298 12499 10301
rect 12801 10298 12867 10301
rect 12433 10296 12867 10298
rect 12433 10240 12438 10296
rect 12494 10240 12806 10296
rect 12862 10240 12867 10296
rect 12433 10238 12867 10240
rect 12433 10235 12499 10238
rect 12801 10235 12867 10238
rect 10593 10162 10659 10165
rect 11789 10162 11855 10165
rect 10593 10160 11855 10162
rect 10593 10104 10598 10160
rect 10654 10104 11794 10160
rect 11850 10104 11855 10160
rect 10593 10102 11855 10104
rect 10593 10099 10659 10102
rect 11789 10099 11855 10102
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 13351 9759 13667 9760
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 8937 9074 9003 9077
rect 11973 9074 12039 9077
rect 12433 9074 12499 9077
rect 8937 9072 12499 9074
rect 8937 9016 8942 9072
rect 8998 9016 11978 9072
rect 12034 9016 12438 9072
rect 12494 9016 12499 9072
rect 8937 9014 12499 9016
rect 8937 9011 9003 9014
rect 11973 9011 12039 9014
rect 12433 9011 12499 9014
rect 15101 8802 15167 8805
rect 15600 8802 16000 8832
rect 15101 8800 16000 8802
rect 15101 8744 15106 8800
rect 15162 8744 16000 8800
rect 15101 8742 16000 8744
rect 15101 8739 15167 8742
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 15600 8712 16000 8742
rect 13351 8671 13667 8672
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15202 8127 15518 8128
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 14917 6898 14983 6901
rect 15600 6898 16000 6928
rect 14917 6896 16000 6898
rect 14917 6840 14922 6896
rect 14978 6840 16000 6896
rect 14917 6838 16000 6840
rect 14917 6835 14983 6838
rect 15600 6808 16000 6838
rect 5717 6762 5783 6765
rect 5901 6762 5967 6765
rect 5717 6760 5967 6762
rect 5717 6704 5722 6760
rect 5778 6704 5906 6760
rect 5962 6704 5967 6760
rect 5717 6702 5967 6704
rect 5717 6699 5783 6702
rect 5901 6699 5967 6702
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 9121 5674 9187 5677
rect 10961 5674 11027 5677
rect 9121 5672 11027 5674
rect 9121 5616 9126 5672
rect 9182 5616 10966 5672
rect 11022 5616 11027 5672
rect 9121 5614 11027 5616
rect 9121 5611 9187 5614
rect 10961 5611 11027 5614
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 8201 5130 8267 5133
rect 10501 5130 10567 5133
rect 8201 5128 10567 5130
rect 8201 5072 8206 5128
rect 8262 5072 10506 5128
rect 10562 5072 10567 5128
rect 8201 5070 10567 5072
rect 8201 5067 8267 5070
rect 10501 5067 10567 5070
rect 15600 4992 16000 5024
rect 15600 4936 15658 4992
rect 15714 4936 16000 4992
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15600 4904 16000 4936
rect 15202 4863 15518 4864
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 14825 3090 14891 3093
rect 15600 3090 16000 3120
rect 14825 3088 16000 3090
rect 14825 3032 14830 3088
rect 14886 3032 16000 3088
rect 14825 3030 16000 3032
rect 14825 3027 14891 3030
rect 15600 3000 16000 3030
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 13813 1186 13879 1189
rect 15600 1186 16000 1216
rect 13813 1184 16000 1186
rect 13813 1128 13818 1184
rect 13874 1128 16000 1184
rect 13813 1126 16000 1128
rect 13813 1123 13879 1126
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 15600 1096 16000 1126
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__o221a_1  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12512 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12696 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _154_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _155_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _157_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11224 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _158_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11684 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11316 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _161_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12788 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _162_
timestamp 1704896540
transform -1 0 13248 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13248 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12880 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12696 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _166_
timestamp 1704896540
transform -1 0 11776 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1704896540
transform 1 0 11500 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13064 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _169_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10396 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 14168 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13800 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _172_
timestamp 1704896540
transform 1 0 12512 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _173_
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _174_
timestamp 1704896540
transform -1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _175_
timestamp 1704896540
transform 1 0 11316 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _176_
timestamp 1704896540
transform -1 0 12604 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _177_
timestamp 1704896540
transform 1 0 11408 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _179_
timestamp 1704896540
transform 1 0 9844 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _180_
timestamp 1704896540
transform 1 0 10304 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1704896540
transform 1 0 10028 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1704896540
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10212 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _185_
timestamp 1704896540
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 1704896540
transform -1 0 8924 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1704896540
transform -1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _188_
timestamp 1704896540
transform 1 0 6256 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _189_
timestamp 1704896540
transform 1 0 7544 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _190_
timestamp 1704896540
transform 1 0 6716 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _191_
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _192_
timestamp 1704896540
transform 1 0 5888 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _193_
timestamp 1704896540
transform 1 0 5612 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _194_
timestamp 1704896540
transform -1 0 5428 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _195_
timestamp 1704896540
transform 1 0 4416 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 1704896540
transform -1 0 6624 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _197_
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _199_
timestamp 1704896540
transform 1 0 6532 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _200_
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _201_
timestamp 1704896540
transform 1 0 4968 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1704896540
transform -1 0 8096 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _203_
timestamp 1704896540
transform 1 0 7728 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _204_
timestamp 1704896540
transform 1 0 7544 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _205_
timestamp 1704896540
transform -1 0 8280 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _206_
timestamp 1704896540
transform 1 0 8280 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _207_
timestamp 1704896540
transform -1 0 9108 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _208_
timestamp 1704896540
transform 1 0 8740 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1704896540
transform -1 0 9476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _210_
timestamp 1704896540
transform -1 0 9384 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp 1704896540
transform -1 0 9752 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _212_
timestamp 1704896540
transform 1 0 8924 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _213_
timestamp 1704896540
transform 1 0 8556 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _214_
timestamp 1704896540
transform -1 0 8280 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _215_
timestamp 1704896540
transform -1 0 7360 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _216_
timestamp 1704896540
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _217_
timestamp 1704896540
transform -1 0 7360 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _218_
timestamp 1704896540
transform -1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _219_
timestamp 1704896540
transform -1 0 8188 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _220_
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _221_
timestamp 1704896540
transform 1 0 6164 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _222_
timestamp 1704896540
transform -1 0 6440 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _223_
timestamp 1704896540
transform 1 0 5060 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _224_
timestamp 1704896540
transform -1 0 6532 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _225_
timestamp 1704896540
transform 1 0 5336 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _226_
timestamp 1704896540
transform -1 0 5336 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1704896540
transform 1 0 3680 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _228_
timestamp 1704896540
transform 1 0 4232 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _229_
timestamp 1704896540
transform -1 0 6440 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _230_
timestamp 1704896540
transform -1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _231_
timestamp 1704896540
transform -1 0 5520 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _232_
timestamp 1704896540
transform -1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _233_
timestamp 1704896540
transform 1 0 6348 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _234_
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1704896540
transform 1 0 14076 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _236_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1704896540
transform -1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _238_
timestamp 1704896540
transform -1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13064 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _240_
timestamp 1704896540
transform -1 0 12604 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 1704896540
transform 1 0 10764 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _242_
timestamp 1704896540
transform 1 0 10304 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _243_
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 1704896540
transform 1 0 10580 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _245_
timestamp 1704896540
transform 1 0 8648 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _246_
timestamp 1704896540
transform 1 0 9200 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 1704896540
transform -1 0 9292 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _248_
timestamp 1704896540
transform 1 0 7820 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _249_
timestamp 1704896540
transform 1 0 8372 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 1704896540
transform 1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _251_
timestamp 1704896540
transform -1 0 7820 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _252_
timestamp 1704896540
transform -1 0 7452 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 1704896540
transform -1 0 6992 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _254_
timestamp 1704896540
transform 1 0 6072 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _255_
timestamp 1704896540
transform -1 0 6532 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 1704896540
transform 1 0 4784 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _257_
timestamp 1704896540
transform -1 0 5612 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _258_
timestamp 1704896540
transform -1 0 5152 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1704896540
transform 1 0 4508 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _260_
timestamp 1704896540
transform -1 0 4968 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _261_
timestamp 1704896540
transform 1 0 4692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _262_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4140 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4876 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _265_
timestamp 1704896540
transform 1 0 6808 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _266_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7268 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _267_
timestamp 1704896540
transform -1 0 9108 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9568 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _269_
timestamp 1704896540
transform 1 0 9568 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _270_
timestamp 1704896540
transform -1 0 8280 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _271_
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _272_
timestamp 1704896540
transform 1 0 8464 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _273_
timestamp 1704896540
transform 1 0 4692 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _274_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3956 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _275_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9016 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _276_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10580 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _277_
timestamp 1704896540
transform 1 0 7084 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _279_
timestamp 1704896540
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1704896540
transform 1 0 11868 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1704896540
transform -1 0 11592 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _282_
timestamp 1704896540
transform -1 0 11868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _283_
timestamp 1704896540
transform -1 0 11500 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _284_
timestamp 1704896540
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _285_
timestamp 1704896540
transform 1 0 11316 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _286_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 13248 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _287_
timestamp 1704896540
transform 1 0 11684 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _288_
timestamp 1704896540
transform 1 0 12512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _289_
timestamp 1704896540
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _290_
timestamp 1704896540
transform -1 0 12512 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _291_
timestamp 1704896540
transform 1 0 12512 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _292_
timestamp 1704896540
transform 1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _293_
timestamp 1704896540
transform 1 0 12972 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1704896540
transform 1 0 12144 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _295_
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _296_
timestamp 1704896540
transform -1 0 12788 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _297_
timestamp 1704896540
transform -1 0 13616 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _298_
timestamp 1704896540
transform -1 0 13984 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _299_
timestamp 1704896540
transform -1 0 13064 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _300_
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _301_
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _302_
timestamp 1704896540
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _304_
timestamp 1704896540
transform 1 0 9384 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _305_
timestamp 1704896540
transform 1 0 9108 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _306_
timestamp 1704896540
transform 1 0 7912 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _307_
timestamp 1704896540
transform 1 0 5980 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _308_
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _309_
timestamp 1704896540
transform -1 0 4140 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _310_
timestamp 1704896540
transform 1 0 3220 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _311_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13340 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _312_
timestamp 1704896540
transform 1 0 13248 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _313_
timestamp 1704896540
transform 1 0 13340 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _314_
timestamp 1704896540
transform 1 0 13340 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _315_
timestamp 1704896540
transform 1 0 13340 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _316_
timestamp 1704896540
transform 1 0 12972 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _317_
timestamp 1704896540
transform -1 0 13340 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _318_
timestamp 1704896540
transform 1 0 13340 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _319_
timestamp 1704896540
transform 1 0 9752 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _320_
timestamp 1704896540
transform -1 0 13248 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _321_
timestamp 1704896540
transform 1 0 9384 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _322_
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _323_
timestamp 1704896540
transform -1 0 8188 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _324_
timestamp 1704896540
transform 1 0 4048 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _325_
timestamp 1704896540
transform 1 0 3404 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _326_
timestamp 1704896540
transform 1 0 3404 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _327_
timestamp 1704896540
transform 1 0 8372 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _328_
timestamp 1704896540
transform -1 0 10580 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _329_
timestamp 1704896540
transform 1 0 9200 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _330_
timestamp 1704896540
transform 1 0 7084 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _331_
timestamp 1704896540
transform 1 0 3956 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _332_
timestamp 1704896540
transform 1 0 3312 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _333_
timestamp 1704896540
transform -1 0 4692 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _334_
timestamp 1704896540
transform 1 0 5796 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _335__12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13616 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _335_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13248 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11040 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1704896540
transform -1 0 7728 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1704896540
transform 1 0 6072 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1704896540
transform 1 0 11592 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1704896540
transform 1 0 11776 0 -1 12512
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1704896540
transform 1 0 9476 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1704896540
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1704896540
transform 1 0 14996 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1704896540
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1704896540
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1704896540
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_106
timestamp 1704896540
transform 1 0 10304 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_118
timestamp 1704896540
transform 1 0 11408 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_130
timestamp 1704896540
transform 1 0 12512 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1704896540
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1704896540
transform 1 0 14996 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_45
timestamp 1704896540
transform 1 0 4692 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_57
timestamp 1704896540
transform 1 0 5796 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_63
timestamp 1704896540
transform 1 0 6348 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_75
timestamp 1704896540
transform 1 0 7452 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_108
timestamp 1704896540
transform 1 0 10488 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_120
timestamp 1704896540
transform 1 0 11592 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_132
timestamp 1704896540
transform 1 0 12696 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1704896540
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_35
timestamp 1704896540
transform 1 0 3772 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1704896540
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_63
timestamp 1704896540
transform 1 0 6348 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_83
timestamp 1704896540
transform 1 0 8188 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_87
timestamp 1704896540
transform 1 0 8556 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_103
timestamp 1704896540
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1704896540
transform 1 0 14996 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_63
timestamp 1704896540
transform 1 0 6348 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_114
timestamp 1704896540
transform 1 0 11040 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_131
timestamp 1704896540
transform 1 0 12604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_138
timestamp 1704896540
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1704896540
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_154
timestamp 1704896540
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1704896540
transform 1 0 4876 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1704896540
transform 1 0 6164 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_67
timestamp 1704896540
transform 1 0 6716 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_75
timestamp 1704896540
transform 1 0 7452 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_80
timestamp 1704896540
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_84
timestamp 1704896540
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_91
timestamp 1704896540
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_97
timestamp 1704896540
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_129
timestamp 1704896540
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_138
timestamp 1704896540
transform 1 0 13248 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_47
timestamp 1704896540
transform 1 0 4876 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_66
timestamp 1704896540
transform 1 0 6624 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_70
timestamp 1704896540
transform 1 0 6992 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_75
timestamp 1704896540
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1704896540
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_97
timestamp 1704896540
transform 1 0 9476 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_116
timestamp 1704896540
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_128
timestamp 1704896540
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_133
timestamp 1704896540
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_152
timestamp 1704896540
transform 1 0 14536 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 1704896540
transform 1 0 4876 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_70
timestamp 1704896540
transform 1 0 6992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_101
timestamp 1704896540
transform 1 0 9844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_107
timestamp 1704896540
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_122
timestamp 1704896540
transform 1 0 11776 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_142
timestamp 1704896540
transform 1 0 13616 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_154
timestamp 1704896540
transform 1 0 14720 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_64
timestamp 1704896540
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_73
timestamp 1704896540
transform 1 0 7268 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_77
timestamp 1704896540
transform 1 0 7636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1704896540
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_109
timestamp 1704896540
transform 1 0 10580 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_150
timestamp 1704896540
transform 1 0 14352 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_83
timestamp 1704896540
transform 1 0 8188 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_97
timestamp 1704896540
transform 1 0 9476 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13156 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_33
timestamp 1704896540
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_74
timestamp 1704896540
transform 1 0 7360 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_109
timestamp 1704896540
transform 1 0 10580 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_132
timestamp 1704896540
transform 1 0 12696 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_149
timestamp 1704896540
transform 1 0 14260 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1704896540
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_46
timestamp 1704896540
transform 1 0 4784 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_74
timestamp 1704896540
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_86
timestamp 1704896540
transform 1 0 8464 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 1704896540
transform 1 0 8832 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_100
timestamp 1704896540
transform 1 0 9752 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12052 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_129
timestamp 1704896540
transform 1 0 12420 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_65
timestamp 1704896540
transform 1 0 6532 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_76
timestamp 1704896540
transform 1 0 7544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_93
timestamp 1704896540
transform 1 0 9108 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_114
timestamp 1704896540
transform 1 0 11040 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_121
timestamp 1704896540
transform 1 0 11684 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_129
timestamp 1704896540
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1704896540
transform 1 0 13064 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_146
timestamp 1704896540
transform 1 0 13984 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_64
timestamp 1704896540
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9108 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1704896540
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_113
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_132
timestamp 1704896540
transform 1 0 12696 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_154
timestamp 1704896540
transform 1 0 14720 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_62
timestamp 1704896540
transform 1 0 6256 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_67
timestamp 1704896540
transform 1 0 6716 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_79
timestamp 1704896540
transform 1 0 7820 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8372 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_100
timestamp 1704896540
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_112
timestamp 1704896540
transform 1 0 10856 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_116
timestamp 1704896540
transform 1 0 11224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1704896540
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 1704896540
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4140 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_47
timestamp 1704896540
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1704896540
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_82
timestamp 1704896540
transform 1 0 8096 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9108 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_97
timestamp 1704896540
transform 1 0 9476 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1704896540
transform 1 0 10580 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_116
timestamp 1704896540
transform 1 0 11224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_127
timestamp 1704896540
transform 1 0 12236 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_37
timestamp 1704896540
transform 1 0 3956 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5428 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_59
timestamp 1704896540
transform 1 0 5980 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 1704896540
transform 1 0 7912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_94
timestamp 1704896540
transform 1 0 9200 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_115
timestamp 1704896540
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_124
timestamp 1704896540
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_129
timestamp 1704896540
transform 1 0 12420 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_134
timestamp 1704896540
transform 1 0 12880 0 1 11424
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_144
timestamp 1704896540
transform 1 0 13800 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_156
timestamp 1704896540
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3036 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1704896540
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_57
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_65
timestamp 1704896540
transform 1 0 6532 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_92
timestamp 1704896540
transform 1 0 9016 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_104
timestamp 1704896540
transform 1 0 10120 0 -1 12512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_142
timestamp 1704896540
transform 1 0 13616 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_154
timestamp 1704896540
transform 1 0 14720 0 -1 12512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_37
timestamp 1704896540
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_49
timestamp 1704896540
transform 1 0 5060 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_65
timestamp 1704896540
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_70
timestamp 1704896540
transform 1 0 6992 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1704896540
transform 1 0 8096 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_91
timestamp 1704896540
transform 1 0 8924 0 1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_102
timestamp 1704896540
transform 1 0 9936 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_114
timestamp 1704896540
transform 1 0 11040 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp 1704896540
transform 1 0 11408 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_132
timestamp 1704896540
transform 1 0 12696 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1704896540
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_148
timestamp 1704896540
transform 1 0 14168 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_156
timestamp 1704896540
transform 1 0 14904 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_15
timestamp 1704896540
transform 1 0 1932 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4140 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_73
timestamp 1704896540
transform 1 0 7268 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_79
timestamp 1704896540
transform 1 0 7820 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_87
timestamp 1704896540
transform 1 0 8556 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_48
timestamp 1704896540
transform 1 0 4968 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_56
timestamp 1704896540
transform 1 0 5704 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_65
timestamp 1704896540
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_75
timestamp 1704896540
transform 1 0 7452 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_93
timestamp 1704896540
transform 1 0 9108 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_105
timestamp 1704896540
transform 1 0 10212 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_114
timestamp 1704896540
transform 1 0 11040 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_118
timestamp 1704896540
transform 1 0 11408 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_144
timestamp 1704896540
transform 1 0 13800 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_150
timestamp 1704896540
transform 1 0 14352 0 1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1704896540
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1704896540
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_78
timestamp 1704896540
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_121
timestamp 1704896540
transform 1 0 11684 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_14
timestamp 1704896540
transform 1 0 1840 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_21
timestamp 1704896540
transform 1 0 2484 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_35
timestamp 1704896540
transform 1 0 3772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_49
timestamp 1704896540
transform 1 0 5060 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_55
timestamp 1704896540
transform 1 0 5612 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_57
timestamp 1704896540
transform 1 0 5796 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_63
timestamp 1704896540
transform 1 0 6348 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_71
timestamp 1704896540
transform 1 0 7084 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1704896540
transform 1 0 7636 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8188 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_91
timestamp 1704896540
transform 1 0 8924 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_95
timestamp 1704896540
transform 1 0 9292 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_101
timestamp 1704896540
transform 1 0 9844 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_105
timestamp 1704896540
transform 1 0 10212 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1704896540
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_113
timestamp 1704896540
transform 1 0 10948 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_119
timestamp 1704896540
transform 1 0 11500 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_127
timestamp 1704896540
transform 1 0 12236 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_133
timestamp 1704896540
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1704896540
transform 1 0 13248 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_148
timestamp 1704896540
transform 1 0 14168 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_156
timestamp 1704896540
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 5704 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 8280 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 14996 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 14536 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 14720 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 14260 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 5428 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12512 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform 1 0 11224 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 9936 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 8648 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 7360 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 6072 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 4784 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 3496 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform -1 0 2484 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 920 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1704896540
transform -1 0 14168 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_27
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_28
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_29
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_30
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_31
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_32
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_33
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_34
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_35
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_36
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_37
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_38
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_39
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_41
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_43
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_45
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_47
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_49
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_51
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_53
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_55
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_59
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_60
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_61
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_62
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_72
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_76
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_77
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_79
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_80
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_81
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_82
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_84
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_85
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_86
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_87
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_89
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_90
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_91
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_94
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_95
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_97
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_99
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_100
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_101
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_102
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_104
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_105
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_106
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_107
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_109
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_110
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_111
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_112
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_114
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_115
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_117
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_119
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_120
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_121
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_122
timestamp 1704896540
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1704896540
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
<< labels >>
rlabel metal2 s 8036 14688 8036 14688 4 VGND
rlabel metal1 s 7958 15232 7958 15232 4 VPWR
rlabel metal2 s 14214 14280 14214 14280 4 _000_
rlabel metal2 s 11914 14246 11914 14246 4 _001_
rlabel metal1 s 10667 14450 10667 14450 4 _002_
rlabel metal1 s 9660 12954 9660 12954 4 _003_
rlabel metal2 s 9062 14246 9062 14246 4 _004_
rlabel metal2 s 6762 14246 6762 14246 4 _005_
rlabel metal1 s 5796 12954 5796 12954 4 _006_
rlabel metal1 s 3920 13362 3920 13362 4 _007_
rlabel metal1 s 4457 14450 4457 14450 4 _008_
rlabel metal1 s 12558 7922 12558 7922 4 _009_
rlabel metal1 s 13478 4658 13478 4658 4 _010_
rlabel metal1 s 13386 5678 13386 5678 4 _011_
rlabel metal1 s 13478 9010 13478 9010 4 _012_
rlabel metal1 s 12190 11050 12190 11050 4 _013_
rlabel metal1 s 13018 10030 13018 10030 4 _014_
rlabel metal2 s 13018 13532 13018 13532 4 _015_
rlabel metal1 s 13248 11322 13248 11322 4 _016_
rlabel metal1 s 10207 6154 10207 6154 4 _017_
rlabel metal1 s 12562 4726 12562 4726 4 _018_
rlabel metal2 s 10074 3366 10074 3366 4 _019_
rlabel metal1 s 8500 5134 8500 5134 4 _020_
rlabel metal1 s 7686 4726 7686 4726 4 _021_
rlabel metal1 s 4416 4250 4416 4250 4 _022_
rlabel metal2 s 4922 5746 4922 5746 4 _023_
rlabel metal1 s 4365 6834 4365 6834 4 _024_
rlabel metal1 s 8494 6902 8494 6902 4 _025_
rlabel metal2 s 9430 8194 9430 8194 4 _026_
rlabel metal1 s 9614 9146 9614 9146 4 _027_
rlabel metal1 s 7206 10166 7206 10166 4 _028_
rlabel metal1 s 5239 8330 5239 8330 4 _029_
rlabel metal1 s 3680 8602 3680 8602 4 _030_
rlabel metal1 s 4692 10234 4692 10234 4 _031_
rlabel metal1 s 6256 10778 6256 10778 4 _032_
rlabel metal2 s 4738 14416 4738 14416 4 _033_
rlabel metal2 s 4554 14212 4554 14212 4 _034_
rlabel metal1 s 4830 11730 4830 11730 4 _035_
rlabel metal1 s 5014 11798 5014 11798 4 _036_
rlabel metal1 s 8970 11628 8970 11628 4 _037_
rlabel metal1 s 8372 12682 8372 12682 4 _038_
rlabel metal2 s 8234 11798 8234 11798 4 _039_
rlabel metal1 s 8648 11322 8648 11322 4 _040_
rlabel metal2 s 9614 11492 9614 11492 4 _041_
rlabel metal1 s 8878 11696 8878 11696 4 _042_
rlabel metal2 s 7498 12614 7498 12614 4 _043_
rlabel metal1 s 9108 11662 9108 11662 4 _044_
rlabel metal1 s 8464 11866 8464 11866 4 _045_
rlabel metal1 s 4508 12342 4508 12342 4 _046_
rlabel metal2 s 8142 12308 8142 12308 4 _047_
rlabel metal1 s 10442 11288 10442 11288 4 _048_
rlabel metal1 s 6486 5270 6486 5270 4 _049_
rlabel metal1 s 9660 10506 9660 10506 4 _050_
rlabel metal3 s 13110 11084 13110 11084 4 _051_
rlabel metal2 s 5474 10812 5474 10812 4 _052_
rlabel metal1 s 11822 8534 11822 8534 4 _053_
rlabel metal1 s 5382 9418 5382 9418 4 _054_
rlabel metal1 s 11500 8330 11500 8330 4 _055_
rlabel metal1 s 10902 11662 10902 11662 4 _056_
rlabel metal1 s 5198 11152 5198 11152 4 _057_
rlabel metal1 s 13110 5338 13110 5338 4 _058_
rlabel metal1 s 4278 9962 4278 9962 4 _059_
rlabel metal1 s 12374 6834 12374 6834 4 _060_
rlabel metal2 s 12282 6970 12282 6970 4 _061_
rlabel metal1 s 12696 5746 12696 5746 4 _062_
rlabel metal1 s 13846 7310 13846 7310 4 _063_
rlabel metal2 s 14030 6800 14030 6800 4 _064_
rlabel metal1 s 12190 11526 12190 11526 4 _065_
rlabel metal2 s 13570 7038 13570 7038 4 _066_
rlabel metal1 s 13018 6698 13018 6698 4 _067_
rlabel metal1 s 13064 9486 13064 9486 4 _068_
rlabel metal2 s 12650 8874 12650 8874 4 _069_
rlabel metal1 s 13156 8602 13156 8602 4 _070_
rlabel metal1 s 12236 8942 12236 8942 4 _071_
rlabel metal1 s 5474 10064 5474 10064 4 _072_
rlabel metal1 s 12098 10166 12098 10166 4 _073_
rlabel metal1 s 12236 9962 12236 9962 4 _074_
rlabel metal1 s 11178 10982 11178 10982 4 _075_
rlabel metal2 s 11546 9792 11546 9792 4 _076_
rlabel metal1 s 11822 11322 11822 11322 4 _077_
rlabel metal2 s 12190 10812 12190 10812 4 _078_
rlabel metal1 s 12558 10540 12558 10540 4 _079_
rlabel metal2 s 12742 12308 12742 12308 4 _080_
rlabel metal1 s 13340 12818 13340 12818 4 _081_
rlabel metal1 s 12512 11866 12512 11866 4 _082_
rlabel metal1 s 11960 12342 11960 12342 4 _083_
rlabel metal1 s 11822 12410 11822 12410 4 _084_
rlabel metal1 s 12604 12954 12604 12954 4 _085_
rlabel metal1 s 12742 11220 12742 11220 4 _086_
rlabel metal2 s 13754 12138 13754 12138 4 _087_
rlabel metal2 s 12834 11356 12834 11356 4 _088_
rlabel metal1 s 10672 6834 10672 6834 4 _089_
rlabel metal1 s 11822 4794 11822 4794 4 _090_
rlabel metal1 s 11730 5236 11730 5236 4 _091_
rlabel metal2 s 10258 4352 10258 4352 4 _092_
rlabel metal1 s 10626 5168 10626 5168 4 _093_
rlabel metal1 s 10320 3978 10320 3978 4 _094_
rlabel metal1 s 10350 2958 10350 2958 4 _095_
rlabel metal1 s 9384 4794 9384 4794 4 _096_
rlabel metal2 s 7130 4658 7130 4658 4 _097_
rlabel metal2 s 8686 5814 8686 5814 4 _098_
rlabel metal1 s 8280 5746 8280 5746 4 _099_
rlabel metal1 s 6808 5542 6808 5542 4 _100_
rlabel metal1 s 7314 5542 7314 5542 4 _101_
rlabel metal2 s 5842 4352 5842 4352 4 _102_
rlabel metal1 s 5290 5168 5290 5168 4 _103_
rlabel metal2 s 5658 4454 5658 4454 4 _104_
rlabel metal1 s 4830 4046 4830 4046 4 _105_
rlabel metal1 s 5382 6800 5382 6800 4 _106_
rlabel metal2 s 5382 5610 5382 5610 4 _107_
rlabel metal1 s 6900 6970 6900 6970 4 _108_
rlabel metal1 s 5474 6869 5474 6869 4 _109_
rlabel metal1 s 7728 6426 7728 6426 4 _110_
rlabel metal1 s 7774 6766 7774 6766 4 _111_
rlabel metal2 s 8970 7990 8970 7990 4 _112_
rlabel metal1 s 9062 10166 9062 10166 4 _113_
rlabel metal1 s 9032 7990 9032 7990 4 _114_
rlabel metal1 s 9200 7922 9200 7922 4 _115_
rlabel metal1 s 9108 9010 9108 9010 4 _116_
rlabel metal2 s 9246 9860 9246 9860 4 _117_
rlabel metal1 s 7866 8806 7866 8806 4 _118_
rlabel metal1 s 7130 8330 7130 8330 4 _119_
rlabel metal1 s 7130 9452 7130 9452 4 _120_
rlabel metal1 s 6979 9146 6979 9146 4 _121_
rlabel metal2 s 6946 9486 6946 9486 4 _122_
rlabel metal2 s 6854 7514 6854 7514 4 _123_
rlabel metal1 s 6624 7514 6624 7514 4 _124_
rlabel metal2 s 5566 9554 5566 9554 4 _125_
rlabel metal2 s 5106 9418 5106 9418 4 _126_
rlabel metal1 s 5106 9996 5106 9996 4 _127_
rlabel metal1 s 5236 9350 5236 9350 4 _128_
rlabel metal2 s 3910 8874 3910 8874 4 _129_
rlabel metal1 s 5152 10098 5152 10098 4 _130_
rlabel metal1 s 5842 10540 5842 10540 4 _131_
rlabel metal2 s 5382 10744 5382 10744 4 _132_
rlabel metal1 s 7314 10642 7314 10642 4 _133_
rlabel metal1 s 6164 10642 6164 10642 4 _134_
rlabel metal2 s 5198 14178 5198 14178 4 _135_
rlabel metal1 s 10074 11152 10074 11152 4 _136_
rlabel metal1 s 10166 6766 10166 6766 4 _137_
rlabel metal1 s 12604 13702 12604 13702 4 _138_
rlabel metal1 s 10442 14008 10442 14008 4 _139_
rlabel metal1 s 10856 14042 10856 14042 4 _140_
rlabel metal2 s 8878 13294 8878 13294 4 _141_
rlabel metal1 s 9154 12818 9154 12818 4 _142_
rlabel metal1 s 8510 14042 8510 14042 4 _143_
rlabel metal1 s 8326 13702 8326 13702 4 _144_
rlabel metal2 s 7590 13702 7590 13702 4 _145_
rlabel metal1 s 7452 13498 7452 13498 4 _146_
rlabel metal1 s 6578 12954 6578 12954 4 _147_
rlabel metal2 s 6486 13260 6486 13260 4 _148_
rlabel metal2 s 4922 13056 4922 13056 4 _149_
rlabel metal1 s 5152 13498 5152 13498 4 _150_
rlabel metal1 s 10994 9520 10994 9520 4 clk
rlabel metal2 s 7682 9792 7682 9792 4 clknet_0_clk
rlabel metal1 s 4048 4658 4048 4658 4 clknet_2_0__leaf_clk
rlabel metal1 s 4094 13396 4094 13396 4 clknet_2_1__leaf_clk
rlabel metal1 s 9614 6222 9614 6222 4 clknet_2_2__leaf_clk
rlabel metal2 s 9154 11696 9154 11696 4 clknet_2_3__leaf_clk
rlabel metal1 s 10182 5066 10182 5066 4 counter\[0\]
rlabel metal2 s 8970 9792 8970 9792 4 counter\[10\]
rlabel metal1 s 8786 11220 8786 11220 4 counter\[11\]
rlabel metal1 s 6900 12274 6900 12274 4 counter\[12\]
rlabel metal1 s 5290 9044 5290 9044 4 counter\[13\]
rlabel metal2 s 4186 12733 4186 12733 4 counter\[14\]
rlabel metal1 s 4922 12682 4922 12682 4 counter\[15\]
rlabel metal1 s 10212 5338 10212 5338 4 counter\[1\]
rlabel metal1 s 10488 4658 10488 4658 4 counter\[2\]
rlabel metal1 s 9982 5270 9982 5270 4 counter\[3\]
rlabel metal1 s 6486 4794 6486 4794 4 counter\[4\]
rlabel metal2 s 6026 4862 6026 4862 4 counter\[5\]
rlabel metal2 s 6026 5950 6026 5950 4 counter\[6\]
rlabel metal1 s 5175 6630 5175 6630 4 counter\[7\]
rlabel metal1 s 9062 9418 9062 9418 4 counter\[8\]
rlabel metal2 s 9890 11424 9890 11424 4 counter\[9\]
rlabel metal1 s 12512 14926 12512 14926 4 data[0]
rlabel metal1 s 11224 14926 11224 14926 4 data[1]
rlabel metal1 s 10028 14926 10028 14926 4 data[2]
rlabel metal2 s 8694 15317 8694 15317 4 data[3]
rlabel metal1 s 7360 14926 7360 14926 4 data[4]
rlabel metal1 s 5980 14926 5980 14926 4 data[5]
rlabel metal2 s 4830 15317 4830 15317 4 data[6]
rlabel metal2 s 3542 15317 3542 15317 4 data[7]
rlabel metal2 s 13202 14756 13202 14756 4 divider\[0\]
rlabel metal2 s 10810 14042 10810 14042 4 divider\[1\]
rlabel metal1 s 10580 13362 10580 13362 4 divider\[2\]
rlabel metal1 s 9292 14586 9292 14586 4 divider\[3\]
rlabel metal1 s 7452 14450 7452 14450 4 divider\[4\]
rlabel metal2 s 6946 11968 6946 11968 4 divider\[5\]
rlabel metal2 s 4830 12954 4830 12954 4 divider\[6\]
rlabel metal2 s 4646 14756 4646 14756 4 divider\[7\]
rlabel metal1 s 2208 14926 2208 14926 4 ext_data
rlabel metal2 s 966 15351 966 15351 4 load_divider
rlabel metal1 s 13846 14926 13846 14926 4 n_rst
rlabel metal1 s 12098 13804 12098 13804 4 net1
rlabel metal1 s 4600 13838 4600 13838 4 net10
rlabel metal2 s 14122 14314 14122 14314 4 net11
rlabel metal1 s 13616 14518 13616 14518 4 net12
rlabel metal2 s 5290 7004 5290 7004 4 net13
rlabel metal2 s 5198 5338 5198 5338 4 net14
rlabel metal1 s 7452 5134 7452 5134 4 net15
rlabel metal1 s 12006 10574 12006 10574 4 net16
rlabel metal1 s 13294 6222 13294 6222 4 net17
rlabel metal1 s 13616 5202 13616 5202 4 net18
rlabel metal1 s 12144 9486 12144 9486 4 net19
rlabel metal2 s 11408 14382 11408 14382 4 net2
rlabel metal2 s 4922 10268 4922 10268 4 net20
rlabel metal1 s 10074 12750 10074 12750 4 net3
rlabel metal1 s 9568 13838 9568 13838 4 net4
rlabel metal2 s 6946 13634 6946 13634 4 net5
rlabel metal1 s 6440 12750 6440 12750 4 net6
rlabel metal1 s 4646 13260 4646 13260 4 net7
rlabel metal1 s 4416 15062 4416 15062 4 net8
rlabel metal1 s 3036 14790 3036 14790 4 net9
rlabel metal3 s 14774 1156 14774 1156 4 r2r_out[0]
rlabel metal3 s 15280 3060 15280 3060 4 r2r_out[1]
rlabel metal1 s 15318 5542 15318 5542 4 r2r_out[2]
rlabel metal2 s 14950 7837 14950 7837 4 r2r_out[3]
rlabel metal1 s 15042 10982 15042 10982 4 r2r_out[4]
rlabel metal1 s 12144 11118 12144 11118 4 r2r_out[5]
rlabel metal1 s 13248 12750 13248 12750 4 r2r_out[6]
rlabel metal1 s 15088 13430 15088 13430 4 r2r_out[7]
rlabel metal1 s 4922 13872 4922 13872 4 rst
flabel metal4 s 15200 496 15520 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 11498 496 11818 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 7796 496 8116 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4094 496 4414 15280 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 13349 496 13669 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 9647 496 9967 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5945 496 6265 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2243 496 2563 15280 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 15014 15600 15070 16000 0 FreeSans 280 90 0 0 clk
port 3 nsew
flabel metal2 s 12438 15600 12494 16000 0 FreeSans 280 90 0 0 data[0]
port 4 nsew
flabel metal2 s 11150 15600 11206 16000 0 FreeSans 280 90 0 0 data[1]
port 5 nsew
flabel metal2 s 9862 15600 9918 16000 0 FreeSans 280 90 0 0 data[2]
port 6 nsew
flabel metal2 s 8574 15600 8630 16000 0 FreeSans 280 90 0 0 data[3]
port 7 nsew
flabel metal2 s 7286 15600 7342 16000 0 FreeSans 280 90 0 0 data[4]
port 8 nsew
flabel metal2 s 5998 15600 6054 16000 0 FreeSans 280 90 0 0 data[5]
port 9 nsew
flabel metal2 s 4710 15600 4766 16000 0 FreeSans 280 90 0 0 data[6]
port 10 nsew
flabel metal2 s 3422 15600 3478 16000 0 FreeSans 280 90 0 0 data[7]
port 11 nsew
flabel metal2 s 2134 15600 2190 16000 0 FreeSans 280 90 0 0 ext_data
port 12 nsew
flabel metal2 s 846 15600 902 16000 0 FreeSans 280 90 0 0 load_divider
port 13 nsew
flabel metal2 s 13726 15600 13782 16000 0 FreeSans 280 90 0 0 n_rst
port 14 nsew
flabel metal3 s 15600 1096 16000 1216 0 FreeSans 600 0 0 0 r2r_out[0]
port 15 nsew
flabel metal3 s 15600 3000 16000 3120 0 FreeSans 600 0 0 0 r2r_out[1]
port 16 nsew
flabel metal3 s 15600 4904 16000 5024 0 FreeSans 600 0 0 0 r2r_out[2]
port 17 nsew
flabel metal3 s 15600 6808 16000 6928 0 FreeSans 600 0 0 0 r2r_out[3]
port 18 nsew
flabel metal3 s 15600 8712 16000 8832 0 FreeSans 600 0 0 0 r2r_out[4]
port 19 nsew
flabel metal3 s 15600 10616 16000 10736 0 FreeSans 600 0 0 0 r2r_out[5]
port 20 nsew
flabel metal3 s 15600 12520 16000 12640 0 FreeSans 600 0 0 0 r2r_out[6]
port 21 nsew
flabel metal3 s 15600 14424 16000 14544 0 FreeSans 600 0 0 0 r2r_out[7]
port 22 nsew
<< properties >>
string FIXED_BBOX 0 0 16000 16000
string GDS_END 874912
string GDS_FILE ../gds/r2r_dac_control.gds
string GDS_START 281042
<< end >>
